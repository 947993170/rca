module rca(
    input wire rstn,
    input wire [2:0] cfg,
    input wire [5:0] clk_cnt_all,
    input wire [7:0] AES_128_out_0,
    input wire [7:0] AES_128_out_1,
    input wire [7:0] AES_128_out_2,
    input wire [7:0] AES_128_out_3,
    input wire [7:0] AES_128_out_4,
    input wire [7:0] AES_128_out_5,
    input wire [7:0] AES_128_out_6,
    input wire [7:0] AES_128_out_7,
    input wire [7:0] AES_128_out_8,
    input wire [7:0] AES_128_out_9,
    input wire [7:0] AES_128_out_10,
    input wire [7:0] AES_128_out_11,
    input wire [7:0] AES_128_out_12,
    input wire [7:0] AES_128_out_13,
    input wire [7:0] AES_192_out_0,
    input wire [7:0] AES_192_out_1,
    input wire [7:0] AES_192_out_2,
    input wire [7:0] AES_192_out_3,
    input wire [7:0] AES_192_out_4,
    input wire [7:0] AES_192_out_5,
    input wire [7:0] AES_192_out_6,
    input wire [7:0] AES_192_out_7,
    input wire [7:0] AES_192_out_8,
    input wire [7:0] AES_192_out_9,
    input wire [7:0] AES_192_out_10,
    input wire [7:0] AES_192_out_11,
    input wire [7:0] AES_192_out_12,
    input wire [7:0] AES_192_out_13,
    input wire [7:0] AES_256_out_0,
    input wire [7:0] AES_256_out_1,
    input wire [7:0] AES_256_out_2,
    input wire [7:0] AES_256_out_3,
    input wire [7:0] AES_256_out_4,
    input wire [7:0] AES_256_out_5,
    input wire [7:0] AES_256_out_6,
    input wire [7:0] AES_256_out_7,
    input wire [7:0] AES_256_out_8,
    input wire [7:0] AES_256_out_9,
    input wire [7:0] AES_256_out_10,
    input wire [7:0] AES_256_out_11,
    input wire [7:0] AES_256_out_12,
    input wire [7:0] AES_256_out_13,
    input wire [7:0] SM4_out_0,
    input wire [7:0] SM4_out_1,
    input wire [7:0] SM4_out_2,
    input wire [7:0] SM4_out_3,
    input wire [7:0] SM4_out_4,
    input wire [7:0] SM4_out_5,
    input wire [7:0] SM4_out_6,
    input wire [7:0] SM4_out_7,
    input wire [7:0] SM4_out_8,
    input wire [7:0] SM4_out_9,
    input wire [7:0] SM4_out_10,
    input wire [7:0] SM4_out_11,
    input wire [7:0] SM4_out_12,
    output reg [31:0] sbox_kout_aes_128_clk_0,
    output reg [127:0] sbox_dout_aes_128_clk_0,
    output reg [127:0] sbox_dout_aes_128_clk_1,
    output reg [31:0] sbox_kout_aes_128_clk_1,
    output reg [31:0] sbox_kout_aes_128_clk_2,
    output reg [127:0] sbox_dout_aes_128_clk_2,
    output reg [127:0] sbox_dout_aes_128_clk_3,
    output reg [31:0] sbox_kout_aes_128_clk_3,
    output reg [31:0] sbox_kout_aes_128_clk_4,
    output reg [127:0] sbox_dout_aes_128_clk_4,
    output reg [127:0] sbox_dout_aes_128_clk_5,
    output reg [31:0] sbox_kout_aes_128_clk_5,
    output reg [31:0] sbox_kout_aes_128_clk_6,
    output reg [127:0] sbox_dout_aes_128_clk_6,
    output reg [127:0] sbox_dout_aes_128_clk_7,
    output reg [31:0] sbox_kout_aes_128_clk_7,
    output reg [31:0] sbox_kout_aes_128_clk_8,
    output reg [127:0] sbox_dout_aes_128_clk_8,
    output reg [127:0] sbox_dout_aes_128_clk_9,
    output reg [31:0] sbox_kout_aes_128_clk_9,
    output reg [31:0] sbox_kout_aes_128_clk_a,
    output reg [127:0] sbox_dout_aes_128_clk_a,
    output reg [127:0] sbox_dout_aes_128_clk_b,
    output reg [31:0] sbox_kout_aes_128_clk_b,
    output reg [31:0] sbox_kout_aes_128_clk_c,
    output reg [127:0] sbox_dout_aes_128_clk_c,
    output reg [127:0] sbox_dout_aes_128_clk_d,
    output reg [31:0] sbox_kout_aes_128_clk_d,
    output reg [31:0] sbox_kout_aes_128_clk_e,
    output reg [127:0] sbox_dout_aes_128_clk_e,
    output reg [127:0] sbox_dout_aes_128_clk_f,
    output reg [31:0] sbox_kout_aes_128_clk_f,
    output reg [31:0] sbox_kout_aes_128_clk_10,
    output reg [127:0] sbox_dout_aes_128_clk_10,
    output reg [127:0] sbox_dout_aes_128_clk_11,
    output reg [31:0] sbox_kout_aes_128_clk_11,
    output reg [31:0] sbox_kout_aes_128_clk_12,
    output reg [127:0] sbox_dout_aes_128_clk_12,
    output reg [127:0] sbox_dout_aes_128_clk_13,
    output reg [31:0] sbox_kout_aes_128_clk_13,
    output reg [31:0] sbox_kout_aes_128_clk_14,
    output reg [127:0] sbox_dout_aes_128_clk_14,
    output reg [127:0] sbox_dout_aes_128_clk_15,
    output reg [31:0] sbox_kout_aes_128_clk_15,
    output reg [31:0] sbox_kout_aes_128_clk_16,
    output reg [127:0] sbox_dout_aes_128_clk_16,
    output reg [127:0] sbox_dout_aes_128_clk_17,
    output reg [31:0] sbox_kout_aes_128_clk_17,
    output reg [31:0] sbox_kout_aes_128_clk_18,
    output reg [127:0] sbox_dout_aes_128_clk_18,
    output reg [127:0] sbox_dout_aes_128_clk_19,
    output reg [31:0] sbox_kout_aes_128_clk_19,
    output reg [31:0] sbox_kout_aes_128_clk_1a,
    output reg [127:0] sbox_dout_aes_128_clk_1a,
    output reg [127:0] sbox_dout_aes_128_clk_1b,
    output reg [31:0] sbox_kout_aes_128_clk_1b,
    output reg [31:0] sbox_kout_aes_128_clk_1c,
    output reg [127:0] sbox_dout_aes_128_clk_1c,
    output reg [127:0] sbox_dout_aes_128_clk_1d,
    output reg [31:0] sbox_kout_aes_128_clk_1d,
    output reg [31:0] sbox_kout_aes_128_clk_1e,
    output reg [127:0] sbox_dout_aes_128_clk_1e,
    output reg [127:0] sbox_dout_aes_128_clk_1f,
    output reg [31:0] sbox_kout_aes_128_clk_1f,
    output reg [31:0] sbox_kout_aes_128_clk_20,
    output reg [127:0] sbox_dout_aes_128_clk_20,
    output reg [127:0] sbox_dout_aes_128_clk_21,
    output reg [31:0] sbox_kout_aes_128_clk_21,
    output reg [31:0] sbox_kout_aes_128_clk_22,
    output reg [127:0] sbox_dout_aes_128_clk_22,
    output reg [127:0] sbox_dout_aes_128_clk_23,
    output reg [31:0] sbox_kout_aes_128_clk_23,
    output reg [31:0] sbox_kout_aes_128_clk_24,
    output reg [127:0] sbox_dout_aes_128_clk_24,
    output reg [127:0] sbox_dout_aes_128_clk_25,
    output reg [31:0] sbox_kout_aes_128_clk_25,
    output reg [31:0] sbox_kout_aes_128_clk_26,
    output reg [127:0] sbox_dout_aes_128_clk_26,
    output reg [127:0] sbox_dout_aes_128_clk_27,
    output reg [31:0] sbox_kout_aes_128_clk_27,
    output reg [31:0] sbox_kout_aes_192_clk_0,
    output reg [127:0] sbox_dout_aes_192_clk_0,
    output reg [127:0] sbox_dout_aes_192_clk_1,
    output reg [31:0] sbox_kout_aes_192_clk_1,
    output reg [127:0] sbox_dout_aes_192_clk_2,
    output reg [127:0] sbox_dout_aes_192_clk_3,
    output reg [31:0] sbox_kout_aes_192_clk_3,
    output reg [127:0] sbox_dout_aes_192_clk_4,
    output reg [31:0] sbox_kout_aes_192_clk_4,
    output reg [31:0] sbox_kout_aes_192_clk_5,
    output reg [127:0] sbox_dout_aes_192_clk_5,
    output reg [127:0] sbox_dout_aes_192_clk_6,
    output reg [31:0] sbox_kout_aes_192_clk_6,
    output reg [127:0] sbox_dout_aes_192_clk_7,
    output reg [127:0] sbox_dout_aes_192_clk_8,
    output reg [31:0] sbox_kout_aes_192_clk_8,
    output reg [127:0] sbox_dout_aes_192_clk_9,
    output reg [31:0] sbox_kout_aes_192_clk_9,
    output reg [31:0] sbox_kout_aes_192_clk_a,
    output reg [127:0] sbox_dout_aes_192_clk_a,
    output reg [127:0] sbox_dout_aes_192_clk_b,
    output reg [31:0] sbox_kout_aes_192_clk_b,
    output reg [127:0] sbox_dout_aes_192_clk_c,
    output reg [127:0] sbox_dout_aes_192_clk_d,
    output reg [31:0] sbox_kout_aes_192_clk_d,
    output reg [127:0] sbox_dout_aes_192_clk_e,
    output reg [31:0] sbox_kout_aes_192_clk_e,
    output reg [31:0] sbox_kout_aes_192_clk_f,
    output reg [127:0] sbox_dout_aes_192_clk_f,
    output reg [127:0] sbox_dout_aes_192_clk_10,
    output reg [31:0] sbox_kout_aes_192_clk_10,
    output reg [127:0] sbox_dout_aes_192_clk_11,
    output reg [127:0] sbox_dout_aes_192_clk_12,
    output reg [31:0] sbox_kout_aes_192_clk_12,
    output reg [127:0] sbox_dout_aes_192_clk_13,
    output reg [31:0] sbox_kout_aes_192_clk_13,
    output reg [31:0] sbox_kout_aes_192_clk_14,
    output reg [127:0] sbox_dout_aes_192_clk_14,
    output reg [127:0] sbox_dout_aes_192_clk_15,
    output reg [31:0] sbox_kout_aes_192_clk_15,
    output reg [127:0] sbox_dout_aes_192_clk_16,
    output reg [127:0] sbox_dout_aes_192_clk_17,
    output reg [31:0] sbox_kout_aes_192_clk_17,
    output reg [127:0] sbox_dout_aes_192_clk_18,
    output reg [31:0] sbox_kout_aes_192_clk_18,
    output reg [31:0] sbox_kout_aes_192_clk_19,
    output reg [127:0] sbox_dout_aes_192_clk_19,
    output reg [127:0] sbox_dout_aes_192_clk_1a,
    output reg [31:0] sbox_kout_aes_192_clk_1a,
    output reg [127:0] sbox_dout_aes_192_clk_1b,
    output reg [127:0] sbox_dout_aes_192_clk_1c,
    output reg [31:0] sbox_kout_aes_192_clk_1c,
    output reg [127:0] sbox_dout_aes_192_clk_1d,
    output reg [31:0] sbox_kout_aes_192_clk_1d,
    output reg [31:0] sbox_kout_aes_192_clk_1e,
    output reg [127:0] sbox_dout_aes_192_clk_1e,
    output reg [127:0] sbox_dout_aes_192_clk_1f,
    output reg [31:0] sbox_kout_aes_192_clk_1f,
    output reg [127:0] sbox_dout_aes_192_clk_20,
    output reg [127:0] sbox_dout_aes_192_clk_21,
    output reg [31:0] sbox_kout_aes_192_clk_21,
    output reg [127:0] sbox_dout_aes_192_clk_22,
    output reg [31:0] sbox_kout_aes_192_clk_22,
    output reg [31:0] sbox_kout_aes_192_clk_23,
    output reg [127:0] sbox_dout_aes_192_clk_23,
    output reg [127:0] sbox_dout_aes_192_clk_24,
    output reg [31:0] sbox_kout_aes_192_clk_24,
    output reg [127:0] sbox_dout_aes_192_clk_25,
    output reg [127:0] sbox_dout_aes_192_clk_26,
    output reg [31:0] sbox_kout_aes_192_clk_26,
    output reg [127:0] sbox_dout_aes_192_clk_27,
    output reg [31:0] sbox_kout_aes_192_clk_27,
    output reg [31:0] sbox_kout_aes_256_clk_0,
    output reg [127:0] sbox_dout_aes_256_clk_0,
    output reg [127:0] sbox_dout_aes_256_clk_1,
    output reg [31:0] sbox_kout_aes_256_clk_1,
    output reg [127:0] sbox_dout_aes_256_clk_2,
    output reg [31:0] sbox_kout_aes_256_clk_2,
    output reg [31:0] sbox_kout_aes_256_clk_3,
    output reg [127:0] sbox_dout_aes_256_clk_3,
    output reg [127:0] sbox_dout_aes_256_clk_4,
    output reg [31:0] sbox_kout_aes_256_clk_4,
    output reg [127:0] sbox_dout_aes_256_clk_5,
    output reg [31:0] sbox_kout_aes_256_clk_5,
    output reg [127:0] sbox_dout_aes_256_clk_6,
    output reg [127:0] sbox_dout_aes_256_clk_7,
    output reg [31:0] sbox_kout_aes_256_clk_7,
    output reg [127:0] sbox_dout_aes_256_clk_8,
    output reg [31:0] sbox_kout_aes_256_clk_8,
    output reg [127:0] sbox_dout_aes_256_clk_9,
    output reg [31:0] sbox_kout_aes_256_clk_a,
    output reg [127:0] sbox_dout_aes_256_clk_a,
    output reg [127:0] sbox_dout_aes_256_clk_b,
    output reg [31:0] sbox_kout_aes_256_clk_b,
    output reg [127:0] sbox_dout_aes_256_clk_c,
    output reg [31:0] sbox_kout_aes_256_clk_c,
    output reg [31:0] sbox_kout_aes_256_clk_d,
    output reg [127:0] sbox_dout_aes_256_clk_d,
    output reg [127:0] sbox_dout_aes_256_clk_e,
    output reg [31:0] sbox_kout_aes_256_clk_e,
    output reg [127:0] sbox_dout_aes_256_clk_f,
    output reg [31:0] sbox_kout_aes_256_clk_f,
    output reg [127:0] sbox_dout_aes_256_clk_10,
    output reg [127:0] sbox_dout_aes_256_clk_11,
    output reg [31:0] sbox_kout_aes_256_clk_11,
    output reg [127:0] sbox_dout_aes_256_clk_12,
    output reg [31:0] sbox_kout_aes_256_clk_12,
    output reg [127:0] sbox_dout_aes_256_clk_13,
    output reg [31:0] sbox_kout_aes_256_clk_14,
    output reg [127:0] sbox_dout_aes_256_clk_14,
    output reg [127:0] sbox_dout_aes_256_clk_15,
    output reg [31:0] sbox_kout_aes_256_clk_15,
    output reg [127:0] sbox_dout_aes_256_clk_16,
    output reg [31:0] sbox_kout_aes_256_clk_16,
    output reg [31:0] sbox_kout_aes_256_clk_17,
    output reg [127:0] sbox_dout_aes_256_clk_17,
    output reg [127:0] sbox_dout_aes_256_clk_18,
    output reg [31:0] sbox_kout_aes_256_clk_18,
    output reg [127:0] sbox_dout_aes_256_clk_19,
    output reg [31:0] sbox_kout_aes_256_clk_19,
    output reg [127:0] sbox_dout_aes_256_clk_1a,
    output reg [127:0] sbox_dout_aes_256_clk_1b,
    output reg [31:0] sbox_kout_aes_256_clk_1b,
    output reg [127:0] sbox_dout_aes_256_clk_1c,
    output reg [31:0] sbox_kout_aes_256_clk_1c,
    output reg [127:0] sbox_dout_aes_256_clk_1d,
    output reg [31:0] sbox_kout_aes_256_clk_1e,
    output reg [127:0] sbox_dout_aes_256_clk_1e,
    output reg [127:0] sbox_dout_aes_256_clk_1f,
    output reg [31:0] sbox_kout_aes_256_clk_1f,
    output reg [127:0] sbox_dout_aes_256_clk_20,
    output reg [31:0] sbox_kout_aes_256_clk_20,
    output reg [31:0] sbox_kout_aes_256_clk_21,
    output reg [127:0] sbox_dout_aes_256_clk_21,
    output reg [127:0] sbox_dout_aes_256_clk_22,
    output reg [31:0] sbox_kout_aes_256_clk_22,
    output reg [127:0] sbox_dout_aes_256_clk_23,
    output reg [31:0] sbox_kout_aes_256_clk_23,
    output reg [127:0] sbox_dout_aes_256_clk_24,
    output reg [127:0] sbox_dout_aes_256_clk_25,
    output reg [31:0] sbox_kout_aes_256_clk_25,
    output reg [127:0] sbox_dout_aes_256_clk_26,
    output reg [31:0] sbox_kout_aes_256_clk_26,
    output reg [127:0] sbox_dout_aes_256_clk_27,
    output reg [31:0] BK_0_round_0,
    output reg [31:0] B_0_round_0,
    output reg [31:0] BK_1_round_1,
    output reg [31:0] B_1_round_1,
    output reg [31:0] BK_0_round_2,
    output reg [31:0] B_0_round_2,
    output reg [31:0] BK_1_round_3,
    output reg [31:0] B_1_round_3,
    output reg [31:0] BK_0_round_4,
    output reg [31:0] B_0_round_4,
    output reg [31:0] BK_1_round_5,
    output reg [31:0] B_1_round_5,
    output reg [31:0] BK_0_round_6,
    output reg [31:0] B_0_round_6,
    output reg [31:0] BK_1_round_7,
    output reg [31:0] B_1_round_7,
    output reg [31:0] BK_0_round_8,
    output reg [31:0] B_0_round_8,
    output reg [31:0] BK_1_round_9,
    output reg [31:0] B_1_round_9,
    output reg [31:0] BK_0_round_10,
    output reg [31:0] B_0_round_10,
    output reg [31:0] BK_1_round_11,
    output reg [31:0] B_1_round_11,
    output reg [31:0] BK_0_round_12,
    output reg [31:0] B_0_round_12,
    output reg [31:0] BK_1_round_13,
    output reg [31:0] B_1_round_13,
    output reg [31:0] BK_0_round_14,
    output reg [31:0] B_0_round_14,
    output reg [31:0] BK_1_round_15,
    output reg [31:0] B_1_round_15,
    output reg [31:0] BK_0_round_16,
    output reg [31:0] B_0_round_16,
    output reg [31:0] BK_1_round_17,
    output reg [31:0] B_1_round_17,
    output reg [31:0] BK_0_round_18,
    output reg [31:0] B_0_round_18,
    output reg [31:0] BK_1_round_19,
    output reg [31:0] B_1_round_19,
    output reg [31:0] BK_0_round_20,
    output reg [31:0] B_0_round_20,
    output reg [31:0] BK_1_round_21,
    output reg [31:0] B_1_round_21,
    output reg [31:0] BK_0_round_22,
    output reg [31:0] B_0_round_22,
    output reg [31:0] BK_1_round_23,
    output reg [31:0] B_1_round_23,
    output reg [31:0] BK_0_round_24,
    output reg [31:0] B_0_round_24,
    output reg [31:0] BK_1_round_25,
    output reg [31:0] B_1_round_25,
    output reg [31:0] BK_0_round_26,
    output reg [31:0] B_0_round_26,
    output reg [31:0] BK_1_round_27,
    output reg [31:0] B_1_round_27,
    output reg [31:0] BK_0_round_28,
    output reg [31:0] B_0_round_28,
    output reg [31:0] BK_1_round_29,
    output reg [31:0] B_1_round_29,
    output reg [31:0] BK_0_round_30,
    output reg [31:0] B_0_round_30,
    output reg [31:0] BK_1_round_31,
    output reg [31:0] B_1_round_31,
    output reg [31:0] BK_0_round_32,
    output reg [31:0] B_0_round_32,
    output reg [31:0] BK_1_round_33,
    output reg [31:0] B_1_round_33,
    output reg [31:0] BK_0_round_34,
    output reg [31:0] B_0_round_34,
    output reg [31:0] BK_1_round_35,
    output reg [31:0] B_1_round_35,
    output reg [31:0] BK_0_round_36,
    output reg [31:0] B_0_round_36,
    output reg [31:0] BK_1_round_37,
    output reg [31:0] B_1_round_37,
    output reg [31:0] BK_0_round_38,
    output reg [31:0] B_0_round_38,
    output reg [31:0] BK_1_round_39,
    output reg [31:0] B_1_round_39,
    output reg [31:0] BK_0_round_40,
    output reg [31:0] B_0_round_40,
    output reg [31:0] BK_1_round_41,
    output reg [31:0] B_1_round_41,
    output reg [31:0] BK_0_round_42,
    output reg [31:0] B_0_round_42,
    output reg [31:0] BK_1_round_43,
    output reg [31:0] B_1_round_43,
    output reg [31:0] BK_0_round_44,
    output reg [31:0] B_0_round_44,
    output reg [31:0] BK_1_round_45,
    output reg [31:0] B_1_round_45,
    output reg [31:0] BK_0_round_46,
    output reg [31:0] B_0_round_46,
    output reg [31:0] BK_1_round_47,
    output reg [31:0] B_1_round_47,
    output reg [31:0] BK_0_round_48,
    output reg [31:0] B_0_round_48,
    output reg [31:0] BK_1_round_49,
    output reg [31:0] B_1_round_49,
    output reg [31:0] BK_0_round_50,
    output reg [31:0] B_0_round_50,
    output reg [31:0] BK_1_round_51,
    output reg [31:0] B_1_round_51,
    output reg [31:0] BK_0_round_52,
    output reg [31:0] B_0_round_52,
    output reg [31:0] BK_1_round_53,
    output reg [31:0] B_1_round_53,
    output reg [31:0] BK_0_round_54,
    output reg [31:0] B_0_round_54,
    output reg [31:0] BK_1_round_55,
    output reg [31:0] B_1_round_55,
    output reg [31:0] BK_0_round_56,
    output reg [31:0] B_0_round_56,
    output reg [31:0] BK_1_round_57,
    output reg [31:0] B_1_round_57,
    output reg [31:0] BK_0_round_58,
    output reg [31:0] B_0_round_58,
    output reg [31:0] BK_1_round_59,
    output reg [31:0] B_1_round_59,
    output reg [31:0] BK_0_round_60,
    output reg [31:0] B_0_round_60,
    output reg [31:0] BK_1_round_61,
    output reg [31:0] B_1_round_61,
    output reg [31:0] BK_0_round_62,
    output reg [31:0] B_0_round_62,
    output reg [31:0] BK_1_round_63,
    output reg [31:0] B_1_round_63,
    output reg [31:0] sbox_kout_aes_192_clk_2,
    output reg [31:0] sbox_kout_aes_192_clk_7,
    output reg [31:0] sbox_kout_aes_192_clk_c,
    output reg [31:0] sbox_kout_aes_192_clk_11,
    output reg [31:0] sbox_kout_aes_192_clk_16,
    output reg [31:0] sbox_kout_aes_192_clk_1b,
    output reg [31:0] sbox_kout_aes_192_clk_20,
    output reg [31:0] sbox_kout_aes_192_clk_25,
    output reg [31:0] sbox_kout_aes_256_clk_6,
    output reg [31:0] sbox_kout_aes_256_clk_9,
    output reg [31:0] sbox_kout_aes_256_clk_10,
    output reg [31:0] sbox_kout_aes_256_clk_13,
    output reg [31:0] sbox_kout_aes_256_clk_1a,
    output reg [31:0] sbox_kout_aes_256_clk_1d,
    output reg [31:0] sbox_kout_aes_256_clk_24,
    output reg [31:0] sbox_kout_aes_256_clk_27
);
always @(*) begin
    sbox_kout_aes_128_clk_0 = 32'h0;
    if (rstn && cfg[2:1] == 2'b00) begin
        case (clk_cnt_all)
            6'h0: begin
                sbox_kout_aes_128_clk_0[31:24] = AES_128_out_0;
                sbox_kout_aes_128_clk_0[23:16] = AES_128_out_1;
                sbox_kout_aes_128_clk_0[15:8]  = AES_128_out_2;
                sbox_kout_aes_128_clk_0[7:0]   = AES_128_out_3;
            end
        endcase
    end
end

always @(*) begin
    sbox_dout_aes_128_clk_0 = 128'h0;
    if (rstn && cfg[2:1] == 2'b00) begin
        case (clk_cnt_all)
            6'h0: begin
                sbox_dout_aes_128_clk_0[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_0[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_0[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_0[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_0[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_0[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_0[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_0[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_0[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_0[55:48]   = AES_128_out_13;
            end
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_1 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_1 = 128'h0;
        case (clk_cnt_all)
            6'h1: begin
                sbox_dout_aes_128_clk_1[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_1[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_1[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_1[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_1[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_1[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_1[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_1[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_1[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_1[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_1 = sbox_dout_aes_128_clk_1;
        endcase
    end else begin
        sbox_dout_aes_128_clk_1 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_1 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_1 = 32'h0;
        case (clk_cnt_all)
            6'h1: begin
                sbox_kout_aes_128_clk_1[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_1[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_1[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_1[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_1 = sbox_kout_aes_128_clk_1;
        endcase
    end else begin
        sbox_kout_aes_128_clk_1 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_2 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_2 = 32'h0;
        case (clk_cnt_all)
            6'h2: begin
                sbox_kout_aes_128_clk_2[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_2[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_2[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_2[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_2 = sbox_kout_aes_128_clk_2;
        endcase
    end else begin
        sbox_kout_aes_128_clk_2 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_2 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_2 = 128'h0;
        case (clk_cnt_all)
            6'h2: begin
                sbox_dout_aes_128_clk_2[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_2[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_2[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_2[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_2[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_2[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_2[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_2[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_2[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_2[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_2 = sbox_dout_aes_128_clk_2;
        endcase
    end else begin
        sbox_dout_aes_128_clk_2 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_3 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_3 = 128'h0;
        case (clk_cnt_all)
            6'h3: begin
                sbox_dout_aes_128_clk_3[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_3[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_3[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_3[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_3[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_3[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_3[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_3[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_3[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_3[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_3 = sbox_dout_aes_128_clk_3;
        endcase
    end else begin
        sbox_dout_aes_128_clk_3 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_3 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_3 = 32'h0;
        case (clk_cnt_all)
            6'h3: begin
                sbox_kout_aes_128_clk_3[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_3[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_3[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_3[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_3 = sbox_kout_aes_128_clk_3;
        endcase
    end else begin
        sbox_kout_aes_128_clk_3 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_4 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_4 = 32'h0;
        case (clk_cnt_all)
            6'h4: begin
                sbox_kout_aes_128_clk_4[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_4[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_4[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_4[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_4 = sbox_kout_aes_128_clk_4;
        endcase
    end else begin
        sbox_kout_aes_128_clk_4 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_4 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_4 = 128'h0;
        case (clk_cnt_all)
            6'h4: begin
                sbox_dout_aes_128_clk_4[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_4[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_4[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_4[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_4[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_4[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_4[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_4[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_4[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_4[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_4 = sbox_dout_aes_128_clk_4;
        endcase
    end else begin
        sbox_dout_aes_128_clk_4 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_5 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_5 = 128'h0;
        case (clk_cnt_all)
            6'h5: begin
                sbox_dout_aes_128_clk_5[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_5[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_5[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_5[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_5[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_5[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_5[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_5[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_5[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_5[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_5 = sbox_dout_aes_128_clk_5;
        endcase
    end else begin
        sbox_dout_aes_128_clk_5 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_5 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_5 = 32'h0;
        case (clk_cnt_all)
            6'h5: begin
                sbox_kout_aes_128_clk_5[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_5[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_5[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_5[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_5 = sbox_kout_aes_128_clk_5;
        endcase
    end else begin
        sbox_kout_aes_128_clk_5 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_6 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_6 = 32'h0;
        case (clk_cnt_all)
            6'h6: begin
                sbox_kout_aes_128_clk_6[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_6[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_6[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_6[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_6 = sbox_kout_aes_128_clk_6;
        endcase
    end else begin
        sbox_kout_aes_128_clk_6 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_6 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_6 = 128'h0;
        case (clk_cnt_all)
            6'h6: begin
                sbox_dout_aes_128_clk_6[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_6[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_6[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_6[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_6[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_6[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_6[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_6[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_6[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_6[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_6 = sbox_dout_aes_128_clk_6;
        endcase
    end else begin
        sbox_dout_aes_128_clk_6 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_7 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_7 = 128'h0;
        case (clk_cnt_all)
            6'h7: begin
                sbox_dout_aes_128_clk_7[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_7[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_7[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_7[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_7[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_7[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_7[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_7[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_7[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_7[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_7 = sbox_dout_aes_128_clk_7;
        endcase
    end else begin
        sbox_dout_aes_128_clk_7 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_7 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_7 = 32'h0;
        case (clk_cnt_all)
            6'h7: begin
                sbox_kout_aes_128_clk_7[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_7[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_7[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_7[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_7 = sbox_kout_aes_128_clk_7;
        endcase
    end else begin
        sbox_kout_aes_128_clk_7 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_8 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_8 = 32'h0;
        case (clk_cnt_all)
            6'h8: begin
                sbox_kout_aes_128_clk_8[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_8[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_8[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_8[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_8 = sbox_kout_aes_128_clk_8;
        endcase
    end else begin
        sbox_kout_aes_128_clk_8 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_8 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_8 = 128'h0;
        case (clk_cnt_all)
            6'h8: begin
                sbox_dout_aes_128_clk_8[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_8[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_8[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_8[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_8[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_8[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_8[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_8[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_8[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_8[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_8 = sbox_dout_aes_128_clk_8;
        endcase
    end else begin
        sbox_dout_aes_128_clk_8 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_9 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_9 = 128'h0;
        case (clk_cnt_all)
            6'h9: begin
                sbox_dout_aes_128_clk_9[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_9[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_9[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_9[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_9[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_9[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_9[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_9[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_9[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_9[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_9 = sbox_dout_aes_128_clk_9;
        endcase
    end else begin
        sbox_dout_aes_128_clk_9 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_9 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_9 = 32'h0;
        case (clk_cnt_all)
            6'h9: begin
                sbox_kout_aes_128_clk_9[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_9[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_9[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_9[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_9 = sbox_kout_aes_128_clk_9;
        endcase
    end else begin
        sbox_kout_aes_128_clk_9 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_a = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_a = 32'h0;
        case (clk_cnt_all)
            6'ha: begin
                sbox_kout_aes_128_clk_a[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_a[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_a[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_a[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_a = sbox_kout_aes_128_clk_a;
        endcase
    end else begin
        sbox_kout_aes_128_clk_a = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_a = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_a = 128'h0;
        case (clk_cnt_all)
            6'ha: begin
                sbox_dout_aes_128_clk_a[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_a[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_a[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_a[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_a[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_a[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_a[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_a[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_a[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_a[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_a = sbox_dout_aes_128_clk_a;
        endcase
    end else begin
        sbox_dout_aes_128_clk_a = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_b = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_b = 128'h0;
        case (clk_cnt_all)
            6'hb: begin
                sbox_dout_aes_128_clk_b[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_b[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_b[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_b[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_b[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_b[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_b[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_b[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_b[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_b[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_b = sbox_dout_aes_128_clk_b;
        endcase
    end else begin
        sbox_dout_aes_128_clk_b = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_b = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_b = 32'h0;
        case (clk_cnt_all)
            6'hb: begin
                sbox_kout_aes_128_clk_b[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_b[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_b[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_b[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_b = sbox_kout_aes_128_clk_b;
        endcase
    end else begin
        sbox_kout_aes_128_clk_b = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_c = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_c = 32'h0;
        case (clk_cnt_all)
            6'hc: begin
                sbox_kout_aes_128_clk_c[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_c[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_c[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_c[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_c = sbox_kout_aes_128_clk_c;
        endcase
    end else begin
        sbox_kout_aes_128_clk_c = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_c = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_c = 128'h0;
        case (clk_cnt_all)
            6'hc: begin
                sbox_dout_aes_128_clk_c[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_c[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_c[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_c[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_c[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_c[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_c[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_c[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_c[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_c[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_c = sbox_dout_aes_128_clk_c;
        endcase
    end else begin
        sbox_dout_aes_128_clk_c = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_d = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_d = 128'h0;
        case (clk_cnt_all)
            6'hd: begin
                sbox_dout_aes_128_clk_d[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_d[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_d[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_d[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_d[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_d[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_d[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_d[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_d[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_d[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_d = sbox_dout_aes_128_clk_d;
        endcase
    end else begin
        sbox_dout_aes_128_clk_d = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_d = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_d = 32'h0;
        case (clk_cnt_all)
            6'hd: begin
                sbox_kout_aes_128_clk_d[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_d[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_d[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_d[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_d = sbox_kout_aes_128_clk_d;
        endcase
    end else begin
        sbox_kout_aes_128_clk_d = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_e = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_e = 32'h0;
        case (clk_cnt_all)
            6'he: begin
                sbox_kout_aes_128_clk_e[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_e[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_e[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_e[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_e = sbox_kout_aes_128_clk_e;
        endcase
    end else begin
        sbox_kout_aes_128_clk_e = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_e = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_e = 128'h0;
        case (clk_cnt_all)
            6'he: begin
                sbox_dout_aes_128_clk_e[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_e[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_e[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_e[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_e[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_e[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_e[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_e[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_e[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_e[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_e = sbox_dout_aes_128_clk_e;
        endcase
    end else begin
        sbox_dout_aes_128_clk_e = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_f = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_f = 128'h0;
        case (clk_cnt_all)
            6'hf: begin
                sbox_dout_aes_128_clk_f[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_f[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_f[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_f[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_f[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_f[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_f[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_f[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_f[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_f[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_f = sbox_dout_aes_128_clk_f;
        endcase
    end else begin
        sbox_dout_aes_128_clk_f = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_f = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_f = 32'h0;
        case (clk_cnt_all)
            6'hf: begin
                sbox_kout_aes_128_clk_f[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_f[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_f[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_f[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_f = sbox_kout_aes_128_clk_f;
        endcase
    end else begin
        sbox_kout_aes_128_clk_f = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_10 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_10 = 32'h0;
        case (clk_cnt_all)
            6'h10: begin
                sbox_kout_aes_128_clk_10[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_10[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_10[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_10[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_10 = sbox_kout_aes_128_clk_10;
        endcase
    end else begin
        sbox_kout_aes_128_clk_10 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_10 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_10 = 128'h0;
        case (clk_cnt_all)
            6'h10: begin
                sbox_dout_aes_128_clk_10[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_10[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_10[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_10[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_10[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_10[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_10[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_10[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_10[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_10[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_10 = sbox_dout_aes_128_clk_10;
        endcase
    end else begin
        sbox_dout_aes_128_clk_10 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_11 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_11 = 128'h0;
        case (clk_cnt_all)
            6'h11: begin
                sbox_dout_aes_128_clk_11[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_11[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_11[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_11[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_11[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_11[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_11[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_11[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_11[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_11[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_11 = sbox_dout_aes_128_clk_11;
        endcase
    end else begin
        sbox_dout_aes_128_clk_11 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_11 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_11 = 32'h0;
        case (clk_cnt_all)
            6'h11: begin
                sbox_kout_aes_128_clk_11[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_11[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_11[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_11[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_11 = sbox_kout_aes_128_clk_11;
        endcase
    end else begin
        sbox_kout_aes_128_clk_11 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_12 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_12 = 32'h0;
        case (clk_cnt_all)
            6'h12: begin
                sbox_kout_aes_128_clk_12[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_12[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_12[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_12[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_12 = sbox_kout_aes_128_clk_12;
        endcase
    end else begin
        sbox_kout_aes_128_clk_12 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_12 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_12 = 128'h0;
        case (clk_cnt_all)
            6'h12: begin
                sbox_dout_aes_128_clk_12[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_12[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_12[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_12[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_12[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_12[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_12[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_12[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_12[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_12[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_12 = sbox_dout_aes_128_clk_12;
        endcase
    end else begin
        sbox_dout_aes_128_clk_12 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_13 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_13 = 128'h0;
        case (clk_cnt_all)
            6'h13: begin
                sbox_dout_aes_128_clk_13[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_13[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_13[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_13[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_13[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_13[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_13[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_13[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_13[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_13[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_13 = sbox_dout_aes_128_clk_13;
        endcase
    end else begin
        sbox_dout_aes_128_clk_13 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_13 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_13 = 32'h0;
        case (clk_cnt_all)
            6'h13: begin
                sbox_kout_aes_128_clk_13[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_13[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_13[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_13[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_13 = sbox_kout_aes_128_clk_13;
        endcase
    end else begin
        sbox_kout_aes_128_clk_13 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_14 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_14 = 32'h0;
        case (clk_cnt_all)
            6'h14: begin
                sbox_kout_aes_128_clk_14[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_14[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_14[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_14[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_14 = sbox_kout_aes_128_clk_14;
        endcase
    end else begin
        sbox_kout_aes_128_clk_14 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_14 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_14 = 128'h0;
        case (clk_cnt_all)
            6'h14: begin
                sbox_dout_aes_128_clk_14[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_14[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_14[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_14[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_14[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_14[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_14[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_14[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_14[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_14[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_14 = sbox_dout_aes_128_clk_14;
        endcase
    end else begin
        sbox_dout_aes_128_clk_14 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_15 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_15 = 128'h0;
        case (clk_cnt_all)
            6'h15: begin
                sbox_dout_aes_128_clk_15[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_15[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_15[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_15[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_15[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_15[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_15[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_15[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_15[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_15[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_15 = sbox_dout_aes_128_clk_15;
        endcase
    end else begin
        sbox_dout_aes_128_clk_15 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_15 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_15 = 32'h0;
        case (clk_cnt_all)
            6'h15: begin
                sbox_kout_aes_128_clk_15[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_15[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_15[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_15[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_15 = sbox_kout_aes_128_clk_15;
        endcase
    end else begin
        sbox_kout_aes_128_clk_15 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_16 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_16 = 32'h0;
        case (clk_cnt_all)
            6'h16: begin
                sbox_kout_aes_128_clk_16[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_16[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_16[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_16[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_16 = sbox_kout_aes_128_clk_16;
        endcase
    end else begin
        sbox_kout_aes_128_clk_16 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_16 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_16 = 128'h0;
        case (clk_cnt_all)
            6'h16: begin
                sbox_dout_aes_128_clk_16[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_16[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_16[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_16[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_16[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_16[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_16[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_16[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_16[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_16[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_16 = sbox_dout_aes_128_clk_16;
        endcase
    end else begin
        sbox_dout_aes_128_clk_16 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_17 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_17 = 128'h0;
        case (clk_cnt_all)
            6'h17: begin
                sbox_dout_aes_128_clk_17[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_17[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_17[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_17[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_17[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_17[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_17[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_17[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_17[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_17[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_17 = sbox_dout_aes_128_clk_17;
        endcase
    end else begin
        sbox_dout_aes_128_clk_17 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_17 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_17 = 32'h0;
        case (clk_cnt_all)
            6'h17: begin
                sbox_kout_aes_128_clk_17[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_17[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_17[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_17[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_17 = sbox_kout_aes_128_clk_17;
        endcase
    end else begin
        sbox_kout_aes_128_clk_17 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_18 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_18 = 32'h0;
        case (clk_cnt_all)
            6'h18: begin
                sbox_kout_aes_128_clk_18[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_18[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_18[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_18[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_18 = sbox_kout_aes_128_clk_18;
        endcase
    end else begin
        sbox_kout_aes_128_clk_18 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_18 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_18 = 128'h0;
        case (clk_cnt_all)
            6'h18: begin
                sbox_dout_aes_128_clk_18[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_18[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_18[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_18[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_18[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_18[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_18[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_18[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_18[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_18[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_18 = sbox_dout_aes_128_clk_18;
        endcase
    end else begin
        sbox_dout_aes_128_clk_18 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_19 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_19 = 128'h0;
        case (clk_cnt_all)
            6'h19: begin
                sbox_dout_aes_128_clk_19[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_19[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_19[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_19[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_19[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_19[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_19[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_19[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_19[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_19[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_19 = sbox_dout_aes_128_clk_19;
        endcase
    end else begin
        sbox_dout_aes_128_clk_19 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_19 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_19 = 32'h0;
        case (clk_cnt_all)
            6'h19: begin
                sbox_kout_aes_128_clk_19[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_19[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_19[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_19[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_19 = sbox_kout_aes_128_clk_19;
        endcase
    end else begin
        sbox_kout_aes_128_clk_19 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_1a = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_1a = 32'h0;
        case (clk_cnt_all)
            6'h1a: begin
                sbox_kout_aes_128_clk_1a[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_1a[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_1a[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_1a[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_1a = sbox_kout_aes_128_clk_1a;
        endcase
    end else begin
        sbox_kout_aes_128_clk_1a = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_1a = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_1a = 128'h0;
        case (clk_cnt_all)
            6'h1a: begin
                sbox_dout_aes_128_clk_1a[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_1a[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_1a[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_1a[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_1a[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_1a[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_1a[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_1a[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_1a[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_1a[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_1a = sbox_dout_aes_128_clk_1a;
        endcase
    end else begin
        sbox_dout_aes_128_clk_1a = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_1b = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_1b = 128'h0;
        case (clk_cnt_all)
            6'h1b: begin
                sbox_dout_aes_128_clk_1b[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_1b[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_1b[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_1b[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_1b[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_1b[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_1b[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_1b[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_1b[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_1b[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_1b = sbox_dout_aes_128_clk_1b;
        endcase
    end else begin
        sbox_dout_aes_128_clk_1b = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_1b = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_1b = 32'h0;
        case (clk_cnt_all)
            6'h1b: begin
                sbox_kout_aes_128_clk_1b[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_1b[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_1b[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_1b[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_1b = sbox_kout_aes_128_clk_1b;
        endcase
    end else begin
        sbox_kout_aes_128_clk_1b = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_1c = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_1c = 32'h0;
        case (clk_cnt_all)
            6'h1c: begin
                sbox_kout_aes_128_clk_1c[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_1c[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_1c[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_1c[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_1c = sbox_kout_aes_128_clk_1c;
        endcase
    end else begin
        sbox_kout_aes_128_clk_1c = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_1c = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_1c = 128'h0;
        case (clk_cnt_all)
            6'h1c: begin
                sbox_dout_aes_128_clk_1c[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_1c[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_1c[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_1c[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_1c[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_1c[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_1c[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_1c[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_1c[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_1c[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_1c = sbox_dout_aes_128_clk_1c;
        endcase
    end else begin
        sbox_dout_aes_128_clk_1c = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_1d = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_1d = 128'h0;
        case (clk_cnt_all)
            6'h1d: begin
                sbox_dout_aes_128_clk_1d[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_1d[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_1d[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_1d[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_1d[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_1d[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_1d[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_1d[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_1d[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_1d[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_1d = sbox_dout_aes_128_clk_1d;
        endcase
    end else begin
        sbox_dout_aes_128_clk_1d = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_1d = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_1d = 32'h0;
        case (clk_cnt_all)
            6'h1d: begin
                sbox_kout_aes_128_clk_1d[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_1d[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_1d[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_1d[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_1d = sbox_kout_aes_128_clk_1d;
        endcase
    end else begin
        sbox_kout_aes_128_clk_1d = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_1e = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_1e = 32'h0;
        case (clk_cnt_all)
            6'h1e: begin
                sbox_kout_aes_128_clk_1e[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_1e[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_1e[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_1e[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_1e = sbox_kout_aes_128_clk_1e;
        endcase
    end else begin
        sbox_kout_aes_128_clk_1e = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_1e = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_1e = 128'h0;
        case (clk_cnt_all)
            6'h1e: begin
                sbox_dout_aes_128_clk_1e[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_1e[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_1e[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_1e[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_1e[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_1e[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_1e[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_1e[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_1e[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_1e[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_1e = sbox_dout_aes_128_clk_1e;
        endcase
    end else begin
        sbox_dout_aes_128_clk_1e = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_1f = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_1f = 128'h0;
        case (clk_cnt_all)
            6'h1f: begin
                sbox_dout_aes_128_clk_1f[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_1f[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_1f[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_1f[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_1f[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_1f[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_1f[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_1f[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_1f[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_1f[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_1f = sbox_dout_aes_128_clk_1f;
        endcase
    end else begin
        sbox_dout_aes_128_clk_1f = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_1f = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_1f = 32'h0;
        case (clk_cnt_all)
            6'h1f: begin
                sbox_kout_aes_128_clk_1f[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_1f[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_1f[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_1f[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_1f = sbox_kout_aes_128_clk_1f;
        endcase
    end else begin
        sbox_kout_aes_128_clk_1f = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_20 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_20 = 32'h0;
        case (clk_cnt_all)
            6'h20: begin
                sbox_kout_aes_128_clk_20[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_20[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_20[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_20[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_20 = sbox_kout_aes_128_clk_20;
        endcase
    end else begin
        sbox_kout_aes_128_clk_20 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_20 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_20 = 128'h0;
        case (clk_cnt_all)
            6'h20: begin
                sbox_dout_aes_128_clk_20[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_20[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_20[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_20[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_20[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_20[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_20[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_20[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_20[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_20[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_20 = sbox_dout_aes_128_clk_20;
        endcase
    end else begin
        sbox_dout_aes_128_clk_20 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_21 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_21 = 128'h0;
        case (clk_cnt_all)
            6'h21: begin
                sbox_dout_aes_128_clk_21[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_21[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_21[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_21[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_21[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_21[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_21[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_21[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_21[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_21[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_21 = sbox_dout_aes_128_clk_21;
        endcase
    end else begin
        sbox_dout_aes_128_clk_21 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_21 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_21 = 32'h0;
        case (clk_cnt_all)
            6'h21: begin
                sbox_kout_aes_128_clk_21[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_21[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_21[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_21[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_21 = sbox_kout_aes_128_clk_21;
        endcase
    end else begin
        sbox_kout_aes_128_clk_21 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_22 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_22 = 32'h0;
        case (clk_cnt_all)
            6'h22: begin
                sbox_kout_aes_128_clk_22[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_22[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_22[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_22[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_22 = sbox_kout_aes_128_clk_22;
        endcase
    end else begin
        sbox_kout_aes_128_clk_22 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_22 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_22 = 128'h0;
        case (clk_cnt_all)
            6'h22: begin
                sbox_dout_aes_128_clk_22[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_22[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_22[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_22[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_22[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_22[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_22[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_22[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_22[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_22[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_22 = sbox_dout_aes_128_clk_22;
        endcase
    end else begin
        sbox_dout_aes_128_clk_22 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_23 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_23 = 128'h0;
        case (clk_cnt_all)
            6'h23: begin
                sbox_dout_aes_128_clk_23[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_23[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_23[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_23[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_23[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_23[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_23[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_23[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_23[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_23[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_23 = sbox_dout_aes_128_clk_23;
        endcase
    end else begin
        sbox_dout_aes_128_clk_23 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_23 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_23 = 32'h0;
        case (clk_cnt_all)
            6'h23: begin
                sbox_kout_aes_128_clk_23[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_23[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_23[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_23[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_23 = sbox_kout_aes_128_clk_23;
        endcase
    end else begin
        sbox_kout_aes_128_clk_23 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_24 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_24 = 32'h0;
        case (clk_cnt_all)
            6'h24: begin
                sbox_kout_aes_128_clk_24[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_24[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_24[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_24[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_24 = sbox_kout_aes_128_clk_24;
        endcase
    end else begin
        sbox_kout_aes_128_clk_24 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_24 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_24 = 128'h0;
        case (clk_cnt_all)
            6'h24: begin
                sbox_dout_aes_128_clk_24[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_24[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_24[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_24[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_24[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_24[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_24[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_24[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_24[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_24[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_24 = sbox_dout_aes_128_clk_24;
        endcase
    end else begin
        sbox_dout_aes_128_clk_24 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_25 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_25 = 128'h0;
        case (clk_cnt_all)
            6'h25: begin
                sbox_dout_aes_128_clk_25[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_25[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_25[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_25[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_25[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_25[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_25[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_25[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_25[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_25[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_25 = sbox_dout_aes_128_clk_25;
        endcase
    end else begin
        sbox_dout_aes_128_clk_25 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_25 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_25 = 32'h0;
        case (clk_cnt_all)
            6'h25: begin
                sbox_kout_aes_128_clk_25[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_25[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_25[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_25[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_25 = sbox_kout_aes_128_clk_25;
        endcase
    end else begin
        sbox_kout_aes_128_clk_25 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_26 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_26 = 32'h0;
        case (clk_cnt_all)
            6'h26: begin
                sbox_kout_aes_128_clk_26[31:24]   = AES_128_out_0;
                sbox_kout_aes_128_clk_26[23:16]   = AES_128_out_1;
                sbox_kout_aes_128_clk_26[15:8]    = AES_128_out_2;
                sbox_kout_aes_128_clk_26[7:0]     = AES_128_out_3;
            end
            default: sbox_kout_aes_128_clk_26 = sbox_kout_aes_128_clk_26;
        endcase
    end else begin
        sbox_kout_aes_128_clk_26 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_26 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_26 = 128'h0;
        case (clk_cnt_all)
            6'h26: begin
                sbox_dout_aes_128_clk_26[127:120] = AES_128_out_4;
                sbox_dout_aes_128_clk_26[119:112] = AES_128_out_5;
                sbox_dout_aes_128_clk_26[111:104] = AES_128_out_6;
                sbox_dout_aes_128_clk_26[103:96]  = AES_128_out_7;
                sbox_dout_aes_128_clk_26[95:88]   = AES_128_out_8;
                sbox_dout_aes_128_clk_26[87:80]   = AES_128_out_9;
                sbox_dout_aes_128_clk_26[79:72]   = AES_128_out_10;
                sbox_dout_aes_128_clk_26[71:64]   = AES_128_out_11;
                sbox_dout_aes_128_clk_26[63:56]   = AES_128_out_12;
                sbox_dout_aes_128_clk_26[55:48]   = AES_128_out_13;
            end
            default: sbox_dout_aes_128_clk_26 = sbox_dout_aes_128_clk_26;
        endcase
    end else begin
        sbox_dout_aes_128_clk_26 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_128_clk_27 = 128'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_dout_aes_128_clk_27 = 128'h0;
        case (clk_cnt_all)
            6'h27: begin
                sbox_dout_aes_128_clk_27[79:72]   = AES_128_out_0;
                sbox_dout_aes_128_clk_27[71:64]   = AES_128_out_1;
                sbox_dout_aes_128_clk_27[63:56]   = AES_128_out_2;
                sbox_dout_aes_128_clk_27[55:48]   = AES_128_out_3;
                sbox_dout_aes_128_clk_27[47:40]   = AES_128_out_4;
                sbox_dout_aes_128_clk_27[39:32]   = AES_128_out_5;
                sbox_dout_aes_128_clk_27[31:24]   = AES_128_out_6;
                sbox_dout_aes_128_clk_27[23:16]   = AES_128_out_7;
                sbox_dout_aes_128_clk_27[15:8]    = AES_128_out_8;
                sbox_dout_aes_128_clk_27[7:0]     = AES_128_out_9;
            end
            default: sbox_dout_aes_128_clk_27 = sbox_dout_aes_128_clk_27;
        endcase
    end else begin
        sbox_dout_aes_128_clk_27 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_128_clk_27 = 32'h0;
    end else if (cfg[2:1] == 2'b00) begin
        sbox_kout_aes_128_clk_27 = 32'h0;
        case (clk_cnt_all)
            6'h27: begin
                sbox_kout_aes_128_clk_27[31:24]   = AES_128_out_10;
                sbox_kout_aes_128_clk_27[23:16]   = AES_128_out_11;
                sbox_kout_aes_128_clk_27[15:8]    = AES_128_out_12;
                sbox_kout_aes_128_clk_27[7:0]     = AES_128_out_13;
            end
            default: sbox_kout_aes_128_clk_27 = sbox_kout_aes_128_clk_27;
        endcase
    end else begin
        sbox_kout_aes_128_clk_27 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_0 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_0 = 32'h0;
        case (clk_cnt_all)
            6'h0: begin
                sbox_kout_aes_192_clk_0[31:24]   = AES_192_out_0;
                sbox_kout_aes_192_clk_0[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_0[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_0[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_0 = sbox_kout_aes_192_clk_0;
        endcase
    end else begin
        sbox_kout_aes_192_clk_0 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_0 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_0 = 128'h0;
        case (clk_cnt_all)
            6'h0: begin
                sbox_dout_aes_192_clk_0[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_0[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_0[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_0[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_0[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_0[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_0[79:72]   = AES_192_out_10;
                sbox_dout_aes_192_clk_0[71:64]   = AES_192_out_11;
                sbox_dout_aes_192_clk_0[63:56]   = AES_192_out_12;
                sbox_dout_aes_192_clk_0[55:48]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_0 = sbox_dout_aes_192_clk_0;
        endcase
    end else begin
        sbox_dout_aes_192_clk_0 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_1 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_1 = 128'h0;
        case (clk_cnt_all)
            6'h1: begin
                sbox_dout_aes_192_clk_1[63:56]   = AES_192_out_0;
                sbox_dout_aes_192_clk_1[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_1[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_1[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_1[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_1[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_1[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_1[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_1[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_1[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_1 = sbox_dout_aes_192_clk_1;
        endcase
    end else begin
        sbox_dout_aes_192_clk_1 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_1 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_1 = 32'h0;
        case (clk_cnt_all)
            6'h1: begin
                sbox_kout_aes_192_clk_1[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_1[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_1[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_1[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_1 = sbox_kout_aes_192_clk_1;
        endcase
    end else begin
        sbox_kout_aes_192_clk_1 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_2 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_2 = 128'h0;
        case (clk_cnt_all)
            6'h2: begin
                sbox_dout_aes_192_clk_2[127:120] = AES_192_out_0;
                sbox_dout_aes_192_clk_2[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_2[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_2[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_2[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_2[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_2[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_2[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_2[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_2[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_2[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_2[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_2[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_2[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_2 = sbox_dout_aes_192_clk_2;
        endcase
    end else begin
        sbox_dout_aes_192_clk_2 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_3 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_3 = 128'h0;
        case (clk_cnt_all)
            6'h3: begin
                sbox_dout_aes_192_clk_3[31:24]   = AES_192_out_0;
                sbox_dout_aes_192_clk_3[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_3[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_3[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_3[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_3[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_3[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_3[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_3[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_3[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_3 = sbox_dout_aes_192_clk_3;
        endcase
    end else begin
        sbox_dout_aes_192_clk_3 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_3 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_3 = 32'h0;
        case (clk_cnt_all)
            6'h3: begin
                sbox_kout_aes_192_clk_3[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_3[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_3[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_3[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_3 = sbox_kout_aes_192_clk_3;
        endcase
    end else begin
        sbox_kout_aes_192_clk_3 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_4 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_4 = 128'h0;
        case (clk_cnt_all)
            6'h4: begin
                sbox_dout_aes_192_clk_4[95:88]   = AES_192_out_0;
                sbox_dout_aes_192_clk_4[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_4[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_4[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_4[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_4[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_4[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_4[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_4[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_4[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_4[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_4[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_4 = sbox_dout_aes_192_clk_4;
        endcase
    end else begin
        sbox_dout_aes_192_clk_4 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_4 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_4 = 32'h0;
        case (clk_cnt_all)
            6'h4: begin
                sbox_kout_aes_192_clk_4[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_4[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_4 = sbox_kout_aes_192_clk_4;
        endcase
    end else begin
        sbox_kout_aes_192_clk_4 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_5 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_5 = 32'h0;
        case (clk_cnt_all)
            6'h5: begin
                sbox_kout_aes_192_clk_5[31:24]   = AES_192_out_0;
                sbox_kout_aes_192_clk_5[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_5[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_5[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_5 = sbox_kout_aes_192_clk_5;
        endcase
    end else begin
        sbox_kout_aes_192_clk_5 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_5 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_5 = 128'h0;
        case (clk_cnt_all)
            6'h5: begin
                sbox_dout_aes_192_clk_5[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_5[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_5[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_5[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_5[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_5[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_5[79:72]   = AES_192_out_10;
                sbox_dout_aes_192_clk_5[71:64]   = AES_192_out_11;
                sbox_dout_aes_192_clk_5[63:56]   = AES_192_out_12;
                sbox_dout_aes_192_clk_5[55:48]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_5 = sbox_dout_aes_192_clk_5;
        endcase
    end else begin
        sbox_dout_aes_192_clk_5 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_6 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_6 = 128'h0;
        case (clk_cnt_all)
            6'h6: begin
                sbox_dout_aes_192_clk_6[63:56]   = AES_192_out_0;
                sbox_dout_aes_192_clk_6[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_6[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_6[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_6[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_6[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_6[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_6[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_6[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_6[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_6 = sbox_dout_aes_192_clk_6;
        endcase
    end else begin
        sbox_dout_aes_192_clk_6 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_6 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_6 = 32'h0;
        case (clk_cnt_all)
            6'h6: begin
                sbox_kout_aes_192_clk_6[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_6[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_6[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_6[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_6 = sbox_kout_aes_192_clk_6;
        endcase
    end else begin
        sbox_kout_aes_192_clk_6 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_7 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_7 = 128'h0;
        case (clk_cnt_all)
            6'h7: begin
                sbox_dout_aes_192_clk_7[127:120] = AES_192_out_0;
                sbox_dout_aes_192_clk_7[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_7[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_7[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_7[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_7[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_7[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_7[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_7[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_7[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_7[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_7[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_7[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_7[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_7 = sbox_dout_aes_192_clk_7;
        endcase
    end else begin
        sbox_dout_aes_192_clk_7 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_8 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_8 = 128'h0;
        case (clk_cnt_all)
            6'h8: begin
                sbox_dout_aes_192_clk_8[31:24]   = AES_192_out_0;
                sbox_dout_aes_192_clk_8[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_8[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_8[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_8[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_8[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_8[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_8[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_8[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_8[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_8 = sbox_dout_aes_192_clk_8;
        endcase
    end else begin
        sbox_dout_aes_192_clk_8 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_8 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_8 = 32'h0;
        case (clk_cnt_all)
            6'h8: begin
                sbox_kout_aes_192_clk_8[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_8[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_8[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_8[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_8 = sbox_kout_aes_192_clk_8;
        endcase
    end else begin
        sbox_kout_aes_192_clk_8 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_9 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_9 = 128'h0;
        case (clk_cnt_all)
            6'h9: begin
                sbox_dout_aes_192_clk_9[95:88]   = AES_192_out_0;
                sbox_dout_aes_192_clk_9[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_9[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_9[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_9[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_9[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_9[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_9[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_9[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_9[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_9[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_9[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_9 = sbox_dout_aes_192_clk_9;
        endcase
    end else begin
        sbox_dout_aes_192_clk_9 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_9 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_9 = 32'h0;
        case (clk_cnt_all)
            6'h9: begin
                sbox_kout_aes_192_clk_9[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_9[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_9 = sbox_kout_aes_192_clk_9;
        endcase
    end else begin
        sbox_kout_aes_192_clk_9 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_a = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_a = 32'h0;
        case (clk_cnt_all)
            6'ha: begin
                sbox_kout_aes_192_clk_a[31:24]   = AES_192_out_0;
                sbox_kout_aes_192_clk_a[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_a[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_a[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_a = sbox_kout_aes_192_clk_a;
        endcase
    end else begin
        sbox_kout_aes_192_clk_a = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_a = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_a = 128'h0;
        case (clk_cnt_all)
            6'ha: begin
                sbox_dout_aes_192_clk_a[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_a[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_a[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_a[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_a[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_a[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_a[79:72]   = AES_192_out_10;
                sbox_dout_aes_192_clk_a[71:64]   = AES_192_out_11;
                sbox_dout_aes_192_clk_a[63:56]   = AES_192_out_12;
                sbox_dout_aes_192_clk_a[55:48]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_a = sbox_dout_aes_192_clk_a;
        endcase
    end else begin
        sbox_dout_aes_192_clk_a = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_b = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_b = 128'h0;
        case (clk_cnt_all)
            6'hb: begin
                sbox_dout_aes_192_clk_b[63:56]   = AES_192_out_0;
                sbox_dout_aes_192_clk_b[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_b[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_b[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_b[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_b[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_b[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_b[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_b[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_b[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_b = sbox_dout_aes_192_clk_b;
        endcase
    end else begin
        sbox_dout_aes_192_clk_b = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_b = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_b = 32'h0;
        case (clk_cnt_all)
            6'hb: begin
                sbox_kout_aes_192_clk_b[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_b[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_b[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_b[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_b = sbox_kout_aes_192_clk_b;
        endcase
    end else begin
        sbox_kout_aes_192_clk_b = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_c = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_c = 128'h0;
        case (clk_cnt_all)
            6'hc: begin
                sbox_dout_aes_192_clk_c[127:120] = AES_192_out_0;
                sbox_dout_aes_192_clk_c[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_c[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_c[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_c[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_c[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_c[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_c[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_c[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_c[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_c[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_c[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_c[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_c[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_c = sbox_dout_aes_192_clk_c;
        endcase
    end else begin
        sbox_dout_aes_192_clk_c = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_d = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_d = 128'h0;
        case (clk_cnt_all)
            6'hd: begin
                sbox_dout_aes_192_clk_d[31:24]   = AES_192_out_0;
                sbox_dout_aes_192_clk_d[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_d[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_d[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_d[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_d[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_d[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_d[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_d[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_d[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_d = sbox_dout_aes_192_clk_d;
        endcase
    end else begin
        sbox_dout_aes_192_clk_d = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_d = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_d = 32'h0;
        case (clk_cnt_all)
            6'hd: begin
                sbox_kout_aes_192_clk_d[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_d[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_d[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_d[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_d = sbox_kout_aes_192_clk_d;
        endcase
    end else begin
        sbox_kout_aes_192_clk_d = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_e = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_e = 128'h0;
        case (clk_cnt_all)
            6'he: begin
                sbox_dout_aes_192_clk_e[95:88]   = AES_192_out_0;
                sbox_dout_aes_192_clk_e[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_e[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_e[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_e[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_e[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_e[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_e[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_e[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_e[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_e[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_e[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_e = sbox_dout_aes_192_clk_e;
        endcase
    end else begin
        sbox_dout_aes_192_clk_e = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_e = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_e = 32'h0;
        case (clk_cnt_all)
            6'he: begin
                sbox_kout_aes_192_clk_e[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_e[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_e = sbox_kout_aes_192_clk_e;
        endcase
    end else begin
        sbox_kout_aes_192_clk_e = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_f = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_f = 32'h0;
        case (clk_cnt_all)
            6'hf: begin
                sbox_kout_aes_192_clk_f[31:24]   = AES_192_out_0;
                sbox_kout_aes_192_clk_f[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_f[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_f[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_f = sbox_kout_aes_192_clk_f;
        endcase
    end else begin
        sbox_kout_aes_192_clk_f = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_f = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_f = 128'h0;
        case (clk_cnt_all)
            6'hf: begin
                sbox_dout_aes_192_clk_f[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_f[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_f[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_f[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_f[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_f[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_f[79:72]   = AES_192_out_10;
                sbox_dout_aes_192_clk_f[71:64]   = AES_192_out_11;
                sbox_dout_aes_192_clk_f[63:56]   = AES_192_out_12;
                sbox_dout_aes_192_clk_f[55:48]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_f = sbox_dout_aes_192_clk_f;
        endcase
    end else begin
        sbox_dout_aes_192_clk_f = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_10 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_10 = 128'h0;
        case (clk_cnt_all)
            6'h10: begin
                sbox_dout_aes_192_clk_10[63:56]   = AES_192_out_0;
                sbox_dout_aes_192_clk_10[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_10[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_10[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_10[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_10[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_10[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_10[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_10[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_10[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_10 = sbox_dout_aes_192_clk_10;
        endcase
    end else begin
        sbox_dout_aes_192_clk_10 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_10 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_10 = 32'h0;
        case (clk_cnt_all)
            6'h10: begin
                sbox_kout_aes_192_clk_10[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_10[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_10[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_10[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_10 = sbox_kout_aes_192_clk_10;
        endcase
    end else begin
        sbox_kout_aes_192_clk_10 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_11 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_11 = 128'h0;
        case (clk_cnt_all)
            6'h11: begin
                sbox_dout_aes_192_clk_11[127:120] = AES_192_out_0;
                sbox_dout_aes_192_clk_11[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_11[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_11[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_11[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_11[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_11[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_11[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_11[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_11[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_11[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_11[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_11[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_11[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_11 = sbox_dout_aes_192_clk_11;
        endcase
    end else begin
        sbox_dout_aes_192_clk_11 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_12 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_12 = 128'h0;
        case (clk_cnt_all)
            6'h12: begin
                sbox_dout_aes_192_clk_12[31:24]   = AES_192_out_0;
                sbox_dout_aes_192_clk_12[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_12[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_12[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_12[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_12[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_12[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_12[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_12[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_12[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_12 = sbox_dout_aes_192_clk_12;
        endcase
    end else begin
        sbox_dout_aes_192_clk_12 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_12 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_12 = 32'h0;
        case (clk_cnt_all)
            6'h12: begin
                sbox_kout_aes_192_clk_12[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_12[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_12[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_12[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_12 = sbox_kout_aes_192_clk_12;
        endcase
    end else begin
        sbox_kout_aes_192_clk_12 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_13 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_13 = 128'h0;
        case (clk_cnt_all)
            6'h13: begin
                sbox_dout_aes_192_clk_13[95:88]   = AES_192_out_0;
                sbox_dout_aes_192_clk_13[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_13[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_13[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_13[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_13[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_13[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_13[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_13[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_13[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_13[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_13[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_13 = sbox_dout_aes_192_clk_13;
        endcase
    end else begin
        sbox_dout_aes_192_clk_13 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_13 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_13 = 32'h0;
        case (clk_cnt_all)
            6'h13: begin
                sbox_kout_aes_192_clk_13[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_13[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_13 = sbox_kout_aes_192_clk_13;
        endcase
    end else begin
        sbox_kout_aes_192_clk_13 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_14 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_14 = 32'h0;
        case (clk_cnt_all)
            6'h14: begin
                sbox_kout_aes_192_clk_14[31:24]    = AES_192_out_0;
                sbox_kout_aes_192_clk_14[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_14[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_14[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_14 = sbox_kout_aes_192_clk_14;
        endcase
    end else begin
        sbox_kout_aes_192_clk_14 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_14 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_14 = 128'h0;
        case (clk_cnt_all)
            6'h14: begin
                sbox_dout_aes_192_clk_14[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_14[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_14[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_14[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_14[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_14[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_14[79:72]   = AES_192_out_10;
                sbox_dout_aes_192_clk_14[71:64]   = AES_192_out_11;
                sbox_dout_aes_192_clk_14[63:56]   = AES_192_out_12;
                sbox_dout_aes_192_clk_14[55:48]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_14 = sbox_dout_aes_192_clk_14;
        endcase
    end else begin
        sbox_dout_aes_192_clk_14 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_15 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_15 = 128'h0;
        case (clk_cnt_all)
            6'h15: begin
                sbox_dout_aes_192_clk_15[63:56]    = AES_192_out_0;
                sbox_dout_aes_192_clk_15[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_15[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_15[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_15[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_15[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_15[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_15[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_15[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_15[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_15 = sbox_dout_aes_192_clk_15;
        endcase
    end else begin
        sbox_dout_aes_192_clk_15 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_15 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_15 = 32'h0;
        case (clk_cnt_all)
            6'h15: begin
                sbox_kout_aes_192_clk_15[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_15[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_15[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_15[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_15 = sbox_kout_aes_192_clk_15;
        endcase
    end else begin
        sbox_kout_aes_192_clk_15 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_16 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_16 = 128'h0;
        case (clk_cnt_all)
            6'h16: begin
                sbox_dout_aes_192_clk_16[127:120]  = AES_192_out_0;
                sbox_dout_aes_192_clk_16[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_16[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_16[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_16[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_16[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_16[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_16[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_16[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_16[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_16[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_16[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_16[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_16[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_16 = sbox_dout_aes_192_clk_16;
        endcase
    end else begin
        sbox_dout_aes_192_clk_16 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_17 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_17 = 128'h0;
        case (clk_cnt_all)
            6'h17: begin
                sbox_dout_aes_192_clk_17[31:24]    = AES_192_out_0;
                sbox_dout_aes_192_clk_17[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_17[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_17[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_17[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_17[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_17[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_17[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_17[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_17[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_17 = sbox_dout_aes_192_clk_17;
        endcase
    end else begin
        sbox_dout_aes_192_clk_17 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_17 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_17 = 32'h0;
        case (clk_cnt_all)
            6'h17: begin
                sbox_kout_aes_192_clk_17[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_17[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_17[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_17[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_17 = sbox_kout_aes_192_clk_17;
        endcase
    end else begin
        sbox_kout_aes_192_clk_17 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_18 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_18 = 128'h0;
        case (clk_cnt_all)
            6'h18: begin
                sbox_dout_aes_192_clk_18[95:88]    = AES_192_out_0;
                sbox_dout_aes_192_clk_18[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_18[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_18[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_18[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_18[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_18[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_18[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_18[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_18[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_18[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_18[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_18 = sbox_dout_aes_192_clk_18;
        endcase
    end else begin
        sbox_dout_aes_192_clk_18 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_18 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_18 = 32'h0;
        case (clk_cnt_all)
            6'h18: begin
                sbox_kout_aes_192_clk_18[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_18[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_18 = sbox_kout_aes_192_clk_18;
        endcase
    end else begin
        sbox_kout_aes_192_clk_18 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_19 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_19 = 32'h0;
        case (clk_cnt_all)
            6'h19: begin
                sbox_kout_aes_192_clk_19[31:24]    = AES_192_out_0;
                sbox_kout_aes_192_clk_19[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_19[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_19[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_19 = sbox_kout_aes_192_clk_19;
        endcase
    end else begin
        sbox_kout_aes_192_clk_19 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_19 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_19 = 128'h0;
        case (clk_cnt_all)
            6'h19: begin
                sbox_dout_aes_192_clk_19[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_19[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_19[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_19[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_19[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_19[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_19[79:72]   = AES_192_out_10;
            end
            default: sbox_dout_aes_192_clk_19 = sbox_dout_aes_192_clk_19;
        endcase
    end else begin
        sbox_dout_aes_192_clk_19 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_1a = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_1a = 128'h0;
        case (clk_cnt_all)
            6'h1a: begin
                sbox_dout_aes_192_clk_1a[63:56]    = AES_192_out_0;
                sbox_dout_aes_192_clk_1a[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_1a[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_1a[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_1a[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_1a[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_1a[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_1a[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_1a[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_1a[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_1a = sbox_dout_aes_192_clk_1a;
        endcase
    end else begin
        sbox_dout_aes_192_clk_1a = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_1a = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_1a = 32'h0;
        case (clk_cnt_all)
            6'h1a: begin
                sbox_kout_aes_192_clk_1a[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_1a[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_1a[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_1a[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_1a = sbox_kout_aes_192_clk_1a;
        endcase
    end else begin
        sbox_kout_aes_192_clk_1a = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_1b = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_1b = 128'h0;
        case (clk_cnt_all)
            6'h1b: begin
                sbox_dout_aes_192_clk_1b[127:120]  = AES_192_out_0;
                sbox_dout_aes_192_clk_1b[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_1b[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_1b[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_1b[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_1b[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_1b[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_1b[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_1b[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_1b[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_1b[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_1b[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_1b[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_1b[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_1b = sbox_dout_aes_192_clk_1b;
        endcase
    end else begin
        sbox_dout_aes_192_clk_1b = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_1c = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_1c = 128'h0;
        case (clk_cnt_all)
            6'h1c: begin
                sbox_dout_aes_192_clk_1c[31:24]    = AES_192_out_0;
                sbox_dout_aes_192_clk_1c[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_1c[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_1c[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_1c[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_1c[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_1c[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_1c[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_1c[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_1c[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_1c = sbox_dout_aes_192_clk_1c;
        endcase
    end else begin
        sbox_dout_aes_192_clk_1c = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_1c = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_1c = 32'h0;
        case (clk_cnt_all)
            6'h1c: begin
                sbox_kout_aes_192_clk_1c[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_1c[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_1c[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_1c[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_1c = sbox_kout_aes_192_clk_1c;
        endcase
    end else begin
        sbox_kout_aes_192_clk_1c = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_1d = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_1d = 128'h0;
        case (clk_cnt_all)
            6'h1d: begin
                sbox_dout_aes_192_clk_1d[95:88]    = AES_192_out_0;
                sbox_dout_aes_192_clk_1d[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_1d[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_1d[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_1d[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_1d[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_1d[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_1d[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_1d[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_1d[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_1d[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_1d[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_1d = sbox_dout_aes_192_clk_1d;
        endcase
    end else begin
        sbox_dout_aes_192_clk_1d = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_1d = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_1d = 32'h0;
        case (clk_cnt_all)
            6'h1d: begin
                sbox_kout_aes_192_clk_1d[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_1d[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_1d = sbox_kout_aes_192_clk_1d;
        endcase
    end else begin
        sbox_kout_aes_192_clk_1d = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_1e = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_1e = 32'h0;
        case (clk_cnt_all)
            6'h1e: begin
                sbox_kout_aes_192_clk_1e[31:24]    = AES_192_out_0;
                sbox_kout_aes_192_clk_1e[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_1e[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_1e[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_1e = sbox_kout_aes_192_clk_1e;
        endcase
    end else begin
        sbox_kout_aes_192_clk_1e = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_1e = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_1e = 128'h0;
        case (clk_cnt_all)
            6'h1e: begin
                sbox_dout_aes_192_clk_1e[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_1e[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_1e[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_1e[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_1e[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_1e[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_1e[79:72]   = AES_192_out_10;
                sbox_dout_aes_192_clk_1e[71:64]   = AES_192_out_11;
                sbox_dout_aes_192_clk_1e[63:56]   = AES_192_out_12;
                sbox_dout_aes_192_clk_1e[55:48]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_1e = sbox_dout_aes_192_clk_1e;
        endcase
    end else begin
        sbox_dout_aes_192_clk_1e = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_1f = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_1f = 128'h0;
        case (clk_cnt_all)
            6'h1f: begin
                sbox_dout_aes_192_clk_1f[63:56]    = AES_192_out_0;
                sbox_dout_aes_192_clk_1f[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_1f[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_1f[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_1f[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_1f[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_1f[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_1f[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_1f[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_1f[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_1f = sbox_dout_aes_192_clk_1f;
        endcase
    end else begin
        sbox_dout_aes_192_clk_1f = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_1f = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_1f = 32'h0;
        case (clk_cnt_all)
            6'h1f: begin
                sbox_kout_aes_192_clk_1f[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_1f[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_1f[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_1f[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_1f = sbox_kout_aes_192_clk_1f;
        endcase
    end else begin
        sbox_kout_aes_192_clk_1f = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_20 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_20 = 128'h0;
        case (clk_cnt_all)
            6'h20: begin
                sbox_dout_aes_192_clk_20[127:120]  = AES_192_out_0;
                sbox_dout_aes_192_clk_20[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_20[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_20[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_20[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_20[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_20[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_20[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_20[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_20[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_20[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_20[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_20[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_20[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_20 = sbox_dout_aes_192_clk_20;
        endcase
    end else begin
        sbox_dout_aes_192_clk_20 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_21 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_21 = 128'h0;
        case (clk_cnt_all)
            6'h21: begin
                sbox_dout_aes_192_clk_21[31:24]    = AES_192_out_0;
                sbox_dout_aes_192_clk_21[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_21[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_21[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_21[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_21[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_21[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_21[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_21[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_21[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_21 = sbox_dout_aes_192_clk_21;
        endcase
    end else begin
        sbox_dout_aes_192_clk_21 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_21 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_21 = 32'h0;
        case (clk_cnt_all)
            6'h21: begin
                sbox_kout_aes_192_clk_21[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_21[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_21[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_21[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_21 = sbox_kout_aes_192_clk_21;
        endcase
    end else begin
        sbox_kout_aes_192_clk_21 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_22 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_22 = 128'h0;
        case (clk_cnt_all)
            6'h22: begin
                sbox_dout_aes_192_clk_22[95:88]    = AES_192_out_0;
                sbox_dout_aes_192_clk_22[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_22[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_22[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_22[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_22[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_22[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_22[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_22[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_22[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_22[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_22[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_22 = sbox_dout_aes_192_clk_22;
        endcase
    end else begin
        sbox_dout_aes_192_clk_22 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_22 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_22 = 32'h0;
        case (clk_cnt_all)
            6'h22: begin
                sbox_kout_aes_192_clk_22[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_22[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_22 = sbox_kout_aes_192_clk_22;
        endcase
    end else begin
        sbox_kout_aes_192_clk_22 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_23 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_23 = 32'h0;
        case (clk_cnt_all)
            6'h23: begin
                sbox_kout_aes_192_clk_23[31:24]    = AES_192_out_0;
                sbox_kout_aes_192_clk_23[23:16]   = AES_192_out_1;
                sbox_kout_aes_192_clk_23[15:8]    = AES_192_out_2;
                sbox_kout_aes_192_clk_23[7:0]     = AES_192_out_3;
            end
            default: sbox_kout_aes_192_clk_23 = sbox_kout_aes_192_clk_23;
        endcase
    end else begin
        sbox_kout_aes_192_clk_23 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_23 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_23 = 128'h0;
        case (clk_cnt_all)
            6'h23: begin
                sbox_dout_aes_192_clk_23[127:120] = AES_192_out_4;
                sbox_dout_aes_192_clk_23[119:112] = AES_192_out_5;
                sbox_dout_aes_192_clk_23[111:104] = AES_192_out_6;
                sbox_dout_aes_192_clk_23[103:96]  = AES_192_out_7;
                sbox_dout_aes_192_clk_23[95:88 ]  = AES_192_out_8;
                sbox_dout_aes_192_clk_23[87:80]   = AES_192_out_9;
                sbox_dout_aes_192_clk_23[79:72]   = AES_192_out_10;
                sbox_dout_aes_192_clk_23[71:64]   = AES_192_out_11;
                sbox_dout_aes_192_clk_23[63:56]   = AES_192_out_12;
                sbox_dout_aes_192_clk_23[55:48]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_23 = sbox_dout_aes_192_clk_23;
        endcase
    end else begin
        sbox_dout_aes_192_clk_23 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_24 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_24 = 128'h0;
        case (clk_cnt_all)
            6'h24: begin
                sbox_dout_aes_192_clk_24[63:56]   = AES_192_out_0;
                sbox_dout_aes_192_clk_24[55:48]   = AES_192_out_1;
                sbox_dout_aes_192_clk_24[47:40]   = AES_192_out_2;
                sbox_dout_aes_192_clk_24[39:32]   = AES_192_out_3;
                sbox_dout_aes_192_clk_24[31:24]   = AES_192_out_4;
                sbox_dout_aes_192_clk_24[23:16]   = AES_192_out_5;
                sbox_dout_aes_192_clk_24[15:8]    = AES_192_out_6;
                sbox_dout_aes_192_clk_24[7:0]     = AES_192_out_7;
                sbox_dout_aes_192_clk_24[127:120] = AES_192_out_12;
                sbox_dout_aes_192_clk_24[119:112] = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_24 = sbox_dout_aes_192_clk_24;
        endcase
    end else begin
        sbox_dout_aes_192_clk_24 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_24 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_24 = 32'h0;
        case (clk_cnt_all)
            6'h24: begin
                sbox_kout_aes_192_clk_24[31:24]   = AES_192_out_8;
                sbox_kout_aes_192_clk_24[23:16]   = AES_192_out_9;
                sbox_kout_aes_192_clk_24[15:8]    = AES_192_out_10;
                sbox_kout_aes_192_clk_24[7:0]     = AES_192_out_11;
            end
            default: sbox_kout_aes_192_clk_24 = sbox_kout_aes_192_clk_24;
        endcase
    end else begin
        sbox_kout_aes_192_clk_24 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_25 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_25 = 128'h0;
        case (clk_cnt_all)
            6'h25: begin
                sbox_dout_aes_192_clk_25[127:120] = AES_192_out_0;
                sbox_dout_aes_192_clk_25[119:112] = AES_192_out_1;
                sbox_dout_aes_192_clk_25[111:104] = AES_192_out_2;
                sbox_dout_aes_192_clk_25[103:96]  = AES_192_out_3;
                sbox_dout_aes_192_clk_25[95:88]   = AES_192_out_4;
                sbox_dout_aes_192_clk_25[87:80]   = AES_192_out_5;
                sbox_dout_aes_192_clk_25[79:72]   = AES_192_out_6;
                sbox_dout_aes_192_clk_25[71:64]   = AES_192_out_7;
                sbox_dout_aes_192_clk_25[63:56]   = AES_192_out_8;
                sbox_dout_aes_192_clk_25[55:48]   = AES_192_out_9;
                sbox_dout_aes_192_clk_25[47:40]   = AES_192_out_10;
                sbox_dout_aes_192_clk_25[39:32]   = AES_192_out_11;
                sbox_dout_aes_192_clk_25[31:24]   = AES_192_out_12;
                sbox_dout_aes_192_clk_25[23:16]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_25 = sbox_dout_aes_192_clk_25;
        endcase
    end else begin
        sbox_dout_aes_192_clk_25 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_26 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_26 = 128'h0;
        case (clk_cnt_all)
            6'h26: begin
                sbox_dout_aes_192_clk_26[31:24]   = AES_192_out_0;
                sbox_dout_aes_192_clk_26[23:16]   = AES_192_out_1;
                sbox_dout_aes_192_clk_26[15:8]    = AES_192_out_2;
                sbox_dout_aes_192_clk_26[7:0]     = AES_192_out_3;
                sbox_dout_aes_192_clk_26[127:120] = AES_192_out_8;
                sbox_dout_aes_192_clk_26[119:112] = AES_192_out_9;
                sbox_dout_aes_192_clk_26[111:104] = AES_192_out_10;
                sbox_dout_aes_192_clk_26[103:96]  = AES_192_out_11;
                sbox_dout_aes_192_clk_26[95:88]   = AES_192_out_12;
                sbox_dout_aes_192_clk_26[87:80]   = AES_192_out_13;
            end
            default: sbox_dout_aes_192_clk_26 = sbox_dout_aes_192_clk_26;
        endcase
    end else begin
        sbox_dout_aes_192_clk_26 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_26 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_26 = 32'h0;
        case (clk_cnt_all)
            6'h26: begin
                sbox_kout_aes_192_clk_26[31:24]   = AES_192_out_4;
                sbox_kout_aes_192_clk_26[23:16]   = AES_192_out_5;
                sbox_kout_aes_192_clk_26[15:8]    = AES_192_out_6;
                sbox_kout_aes_192_clk_26[7:0]     = AES_192_out_7;
            end
            default: sbox_kout_aes_192_clk_26 = sbox_kout_aes_192_clk_26;
        endcase
    end else begin
        sbox_kout_aes_192_clk_26 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_192_clk_27 = 128'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_dout_aes_192_clk_27 = 128'h0;
        case (clk_cnt_all)
            6'h27: begin
                sbox_dout_aes_192_clk_27[95:88]   = AES_192_out_0;
                sbox_dout_aes_192_clk_27[87:80]   = AES_192_out_1;
                sbox_dout_aes_192_clk_27[79:72]   = AES_192_out_2;
                sbox_dout_aes_192_clk_27[71:64]   = AES_192_out_3;
                sbox_dout_aes_192_clk_27[63:56]   = AES_192_out_4;
                sbox_dout_aes_192_clk_27[55:48]   = AES_192_out_5;
                sbox_dout_aes_192_clk_27[47:40]   = AES_192_out_6;
                sbox_dout_aes_192_clk_27[39:32]   = AES_192_out_7;
                sbox_dout_aes_192_clk_27[31:24]   = AES_192_out_8;
                sbox_dout_aes_192_clk_27[23:16]   = AES_192_out_9;
                sbox_dout_aes_192_clk_27[15:8]    = AES_192_out_10;
                sbox_dout_aes_192_clk_27[7:0]     = AES_192_out_11;
            end
            default: sbox_dout_aes_192_clk_27 = sbox_dout_aes_192_clk_27;
        endcase
    end else begin
        sbox_dout_aes_192_clk_27 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_27 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_27 = 32'h0;
        case (clk_cnt_all)
            6'h27: begin
                sbox_kout_aes_192_clk_27[31:24]   = AES_192_out_12;
                sbox_kout_aes_192_clk_27[23:16]   = AES_192_out_13;
            end
            default: sbox_kout_aes_192_clk_27 = sbox_kout_aes_192_clk_27;
        endcase
    end else begin
        sbox_kout_aes_192_clk_27 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_0 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_0 = 32'h0;
        case (clk_cnt_all)
            6'h0: begin
                sbox_kout_aes_256_clk_0[31:24]   = AES_256_out_0;
                sbox_kout_aes_256_clk_0[23:16]   = AES_256_out_1;
                sbox_kout_aes_256_clk_0[15:8 ]   = AES_256_out_2;
                sbox_kout_aes_256_clk_0[7:0]     = AES_256_out_3;
            end
            default: sbox_kout_aes_256_clk_0 = sbox_kout_aes_256_clk_0;
        endcase
    end else begin
        sbox_kout_aes_256_clk_0 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_0 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_0 = 128'h0;
        case (clk_cnt_all)
            6'h0: begin
                sbox_dout_aes_256_clk_0[127:120] = AES_256_out_4;
                sbox_dout_aes_256_clk_0[119:112] = AES_256_out_5;
                sbox_dout_aes_256_clk_0[111:104] = AES_256_out_6;
                sbox_dout_aes_256_clk_0[103:96]  = AES_256_out_7;
                sbox_dout_aes_256_clk_0[95:88]   = AES_256_out_8;
                sbox_dout_aes_256_clk_0[87:80]   = AES_256_out_9;
                sbox_dout_aes_256_clk_0[79:72]   = AES_256_out_10;
                sbox_dout_aes_256_clk_0[71:64]   = AES_256_out_11;
                sbox_dout_aes_256_clk_0[63:56]   = AES_256_out_12;
                sbox_dout_aes_256_clk_0[55:48]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_0 = sbox_dout_aes_256_clk_0;
        endcase
    end else begin
        sbox_dout_aes_256_clk_0 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_1 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_1 = 128'h0;
        case (clk_cnt_all)
            6'h1: begin
                sbox_dout_aes_256_clk_1[47:40]   = AES_256_out_0;
                sbox_dout_aes_256_clk_1[39:32]   = AES_256_out_1;
                sbox_dout_aes_256_clk_1[31:24]   = AES_256_out_2;
                sbox_dout_aes_256_clk_1[23:16]   = AES_256_out_3;
                sbox_dout_aes_256_clk_1[15:8]    = AES_256_out_4;
                sbox_dout_aes_256_clk_1[7:0]     = AES_256_out_5;
                sbox_dout_aes_256_clk_1[127:120] = AES_256_out_10;
                sbox_dout_aes_256_clk_1[119:112] = AES_256_out_11;
                sbox_dout_aes_256_clk_1[111:104] = AES_256_out_12;
                sbox_dout_aes_256_clk_1[103:96]  = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_1 = sbox_dout_aes_256_clk_1;
        endcase
    end else begin
        sbox_dout_aes_256_clk_1 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_1 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_1 = 32'h0;
        case (clk_cnt_all)
            6'h1: begin
                sbox_kout_aes_256_clk_1[31:24]   = AES_256_out_6;
                sbox_kout_aes_256_clk_1[23:16]   = AES_256_out_7;
                sbox_kout_aes_256_clk_1[15:8]    = AES_256_out_8;
                sbox_kout_aes_256_clk_1[7:0]     = AES_256_out_9;
            end
            default: sbox_kout_aes_256_clk_1 = sbox_kout_aes_256_clk_1;
        endcase
    end else begin
        sbox_kout_aes_256_clk_1 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_2 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_2 = 128'h0;
        case (clk_cnt_all)
            6'h2: begin
                sbox_dout_aes_256_clk_2[95:88]   = AES_256_out_0;
                sbox_dout_aes_256_clk_2[87:80]   = AES_256_out_1;
                sbox_dout_aes_256_clk_2[79:72]   = AES_256_out_2;
                sbox_dout_aes_256_clk_2[71:64]   = AES_256_out_3;
                sbox_dout_aes_256_clk_2[63:56]   = AES_256_out_4;
                sbox_dout_aes_256_clk_2[55:48]   = AES_256_out_5;
                sbox_dout_aes_256_clk_2[47:40]   = AES_256_out_6;
                sbox_dout_aes_256_clk_2[39:32]   = AES_256_out_7;
                sbox_dout_aes_256_clk_2[31:24]   = AES_256_out_8;
                sbox_dout_aes_256_clk_2[23:16]   = AES_256_out_9;
                sbox_dout_aes_256_clk_2[15:8]    = AES_256_out_10;
                sbox_dout_aes_256_clk_2[7:0]     = AES_256_out_11;
            end
            default: sbox_dout_aes_256_clk_2 = sbox_dout_aes_256_clk_2;
        endcase
    end else begin
        sbox_dout_aes_256_clk_2 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_2 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_2 = 32'h0;
        case (clk_cnt_all)
            6'h2: begin
                sbox_kout_aes_256_clk_2[31:24]   = AES_256_out_12;
                sbox_kout_aes_256_clk_2[23:16]   = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_2 = sbox_kout_aes_256_clk_2;
        endcase
    end else begin
        sbox_kout_aes_256_clk_2 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_3 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_3 = 32'h0;
        case (clk_cnt_all)
            6'h3: begin
                sbox_kout_aes_256_clk_3[15:8]    = AES_256_out_0;
                sbox_kout_aes_256_clk_3[7:0]     = AES_256_out_1;
            end
            default: sbox_kout_aes_256_clk_3 = sbox_kout_aes_256_clk_3;
        endcase
    end else begin
        sbox_kout_aes_256_clk_3 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_3 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_3 = 128'h0;
        case (clk_cnt_all)
            6'h3: begin
                sbox_dout_aes_256_clk_3[127:120] = AES_256_out_2;
                sbox_dout_aes_256_clk_3[119:112] = AES_256_out_3;
                sbox_dout_aes_256_clk_3[111:104] = AES_256_out_4;
                sbox_dout_aes_256_clk_3[103:96]  = AES_256_out_5;
                sbox_dout_aes_256_clk_3[95:88]   = AES_256_out_6;
                sbox_dout_aes_256_clk_3[87:80]   = AES_256_out_7;
                sbox_dout_aes_256_clk_3[79:72]   = AES_256_out_8;
                sbox_dout_aes_256_clk_3[71:64]   = AES_256_out_9;
                sbox_dout_aes_256_clk_3[63:56]   = AES_256_out_10;
                sbox_dout_aes_256_clk_3[55:48]   = AES_256_out_11;
                sbox_dout_aes_256_clk_3[47:40]   = AES_256_out_12;
                sbox_dout_aes_256_clk_3[39:32]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_3 = sbox_dout_aes_256_clk_3;
        endcase
    end else begin
        sbox_dout_aes_256_clk_3 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_4 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_4 = 128'h0;
        case (clk_cnt_all)
            6'h4: begin
                sbox_dout_aes_256_clk_4[31:24]   = AES_256_out_0;
                sbox_dout_aes_256_clk_4[23:16]   = AES_256_out_1;
                sbox_dout_aes_256_clk_4[15:8]    = AES_256_out_2;
                sbox_dout_aes_256_clk_4[7:0]     = AES_256_out_3;
                sbox_dout_aes_256_clk_4[127:120] = AES_256_out_8;
                sbox_dout_aes_256_clk_4[119:112] = AES_256_out_9;
                sbox_dout_aes_256_clk_4[111:104] = AES_256_out_10;
                sbox_dout_aes_256_clk_4[103:96]  = AES_256_out_11;
                sbox_dout_aes_256_clk_4[95:88]   = AES_256_out_12;
                sbox_dout_aes_256_clk_4[87:80]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_4 = sbox_dout_aes_256_clk_4;
        endcase
    end else begin
        sbox_dout_aes_256_clk_4 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_4 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_4 = 32'h0;
        case (clk_cnt_all)
            6'h4: begin
                sbox_kout_aes_256_clk_4[31:24]   = AES_256_out_4;
                sbox_kout_aes_256_clk_4[23:16]   = AES_256_out_5;
                sbox_kout_aes_256_clk_4[15:8]    = AES_256_out_6;
                sbox_kout_aes_256_clk_4[7:0]     = AES_256_out_7;
            end
            default: sbox_kout_aes_256_clk_4 = sbox_kout_aes_256_clk_4;
        endcase
    end else begin
        sbox_kout_aes_256_clk_4 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_5 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_5 = 128'h0;
        case (clk_cnt_all)
            6'h5: begin
                sbox_dout_aes_256_clk_5[79:72]   = AES_256_out_0;
                sbox_dout_aes_256_clk_5[71:64]   = AES_256_out_1;
                sbox_dout_aes_256_clk_5[63:56]   = AES_256_out_2;
                sbox_dout_aes_256_clk_5[55:48]   = AES_256_out_3;
                sbox_dout_aes_256_clk_5[47:40]   = AES_256_out_4;
                sbox_dout_aes_256_clk_5[39:32]   = AES_256_out_5;
                sbox_dout_aes_256_clk_5[31:24]   = AES_256_out_6;
                sbox_dout_aes_256_clk_5[23:16]   = AES_256_out_7;
                sbox_dout_aes_256_clk_5[15:8]    = AES_256_out_8;
                sbox_dout_aes_256_clk_5[7:0]     = AES_256_out_9;
            end
            default: sbox_dout_aes_256_clk_5 = sbox_dout_aes_256_clk_5;
        endcase
    end else begin
        sbox_dout_aes_256_clk_5 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_5 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_5 = 32'h0;
        case (clk_cnt_all)
            6'h5: begin
                sbox_kout_aes_256_clk_5[31:24]   = AES_256_out_10;
                sbox_kout_aes_256_clk_5[23:16]   = AES_256_out_11;
                sbox_kout_aes_256_clk_5[15:8]    = AES_256_out_12;
                sbox_kout_aes_256_clk_5[7:0]     = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_5 = sbox_kout_aes_256_clk_5;
        endcase
    end else begin
        sbox_kout_aes_256_clk_5 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_6 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_6 = 128'h0;
        case (clk_cnt_all)
            6'h6: begin
                sbox_dout_aes_256_clk_6[127:120] = AES_256_out_0;
                sbox_dout_aes_256_clk_6[119:112] = AES_256_out_1;
                sbox_dout_aes_256_clk_6[111:104] = AES_256_out_2;
                sbox_dout_aes_256_clk_6[103:96]  = AES_256_out_3;
                sbox_dout_aes_256_clk_6[95:88]   = AES_256_out_4;
                sbox_dout_aes_256_clk_6[87:80]   = AES_256_out_5;
                sbox_dout_aes_256_clk_6[79:72]   = AES_256_out_6;
                sbox_dout_aes_256_clk_6[71:64]   = AES_256_out_7;
                sbox_dout_aes_256_clk_6[63:56]   = AES_256_out_8;
                sbox_dout_aes_256_clk_6[55:48]   = AES_256_out_9;
                sbox_dout_aes_256_clk_6[47:40]   = AES_256_out_10;
                sbox_dout_aes_256_clk_6[39:32]   = AES_256_out_11;
                sbox_dout_aes_256_clk_6[31:24]   = AES_256_out_12;
                sbox_dout_aes_256_clk_6[23:16]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_6 = sbox_dout_aes_256_clk_6;
        endcase
    end else begin
        sbox_dout_aes_256_clk_6 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_7 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_7 = 128'h0;
        case (clk_cnt_all)
            6'h7: begin
                sbox_dout_aes_256_clk_7[15:8]    = AES_256_out_0;
                sbox_dout_aes_256_clk_7[7:0]     = AES_256_out_1;
                sbox_dout_aes_256_clk_7[127:120] = AES_256_out_6;
                sbox_dout_aes_256_clk_7[119:112] = AES_256_out_7;
                sbox_dout_aes_256_clk_7[111:104] = AES_256_out_8;
                sbox_dout_aes_256_clk_7[103:96]  = AES_256_out_9;
                sbox_dout_aes_256_clk_7[95:88]   = AES_256_out_10;
                sbox_dout_aes_256_clk_7[87:80]   = AES_256_out_11;
                sbox_dout_aes_256_clk_7[79:72]   = AES_256_out_12;
                sbox_dout_aes_256_clk_7[71:64]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_7 = sbox_dout_aes_256_clk_7;
        endcase
    end else begin
        sbox_dout_aes_256_clk_7 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_7 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_7 = 32'h0;
        case (clk_cnt_all)
            6'h7: begin
                sbox_kout_aes_256_clk_7[31:24]   = AES_256_out_2;
                sbox_kout_aes_256_clk_7[23:16]   = AES_256_out_3;
                sbox_kout_aes_256_clk_7[15:8]    = AES_256_out_4;
                sbox_kout_aes_256_clk_7[7:0]     = AES_256_out_5;
            end
            default: sbox_kout_aes_256_clk_7 = sbox_kout_aes_256_clk_7;
        endcase
    end else begin
        sbox_kout_aes_256_clk_7 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_8 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_8 = 128'h0;
        case (clk_cnt_all)
            6'h8: begin
                sbox_dout_aes_256_clk_8[63:56]   = AES_256_out_0;
                sbox_dout_aes_256_clk_8[55:48]   = AES_256_out_1;
                sbox_dout_aes_256_clk_8[47:40]   = AES_256_out_2;
                sbox_dout_aes_256_clk_8[39:32]   = AES_256_out_3;
                sbox_dout_aes_256_clk_8[31:24]   = AES_256_out_4;
                sbox_dout_aes_256_clk_8[23:16]   = AES_256_out_5;
                sbox_dout_aes_256_clk_8[15:8]    = AES_256_out_6;
                sbox_dout_aes_256_clk_8[7:0]     = AES_256_out_7;
                sbox_dout_aes_256_clk_8[127:120] = AES_256_out_12;
                sbox_dout_aes_256_clk_8[119:112] = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_8 = sbox_dout_aes_256_clk_8;
        endcase
    end else begin
        sbox_dout_aes_256_clk_8 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_8 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_8 = 32'h0;
        case (clk_cnt_all)
            6'h8: begin
                sbox_kout_aes_256_clk_8[31:24]   = AES_256_out_8;
                sbox_kout_aes_256_clk_8[23:16]   = AES_256_out_9;
                sbox_kout_aes_256_clk_8[15:8]    = AES_256_out_10;
                sbox_kout_aes_256_clk_8[7:0]     = AES_256_out_11;
            end
            default: sbox_kout_aes_256_clk_8 = sbox_kout_aes_256_clk_8;
        endcase
    end else begin
        sbox_kout_aes_256_clk_8 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_9 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_9 = 128'h0;
        case (clk_cnt_all)
            6'h9: begin
                sbox_dout_aes_256_clk_9[111:104] = AES_256_out_0;
                sbox_dout_aes_256_clk_9[103:96]  = AES_256_out_1;
                sbox_dout_aes_256_clk_9[95:88]   = AES_256_out_2;
                sbox_dout_aes_256_clk_9[87:80]   = AES_256_out_3;
                sbox_dout_aes_256_clk_9[79:72]   = AES_256_out_4;
                sbox_dout_aes_256_clk_9[71:64]   = AES_256_out_5;
                sbox_dout_aes_256_clk_9[63:56]   = AES_256_out_6;
                sbox_dout_aes_256_clk_9[55:48]   = AES_256_out_7;
                sbox_dout_aes_256_clk_9[47:40]   = AES_256_out_8;
                sbox_dout_aes_256_clk_9[39:32]   = AES_256_out_9;
                sbox_dout_aes_256_clk_9[31:24]   = AES_256_out_10;
                sbox_dout_aes_256_clk_9[23:16]   = AES_256_out_11;
                sbox_dout_aes_256_clk_9[15:8]    = AES_256_out_12;
                sbox_dout_aes_256_clk_9[7:0]     = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_9 = sbox_dout_aes_256_clk_9;
        endcase
    end else begin
        sbox_dout_aes_256_clk_9 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_a = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_a = 32'h0;
        case (clk_cnt_all)
            6'ha: begin
                sbox_kout_aes_256_clk_a[31:24]   = AES_256_out_0;
                sbox_kout_aes_256_clk_a[23:16]   = AES_256_out_1;
                sbox_kout_aes_256_clk_a[15:8 ]   = AES_256_out_2;
                sbox_kout_aes_256_clk_a[7:0]     = AES_256_out_3;
            end
            default: sbox_kout_aes_256_clk_a = sbox_kout_aes_256_clk_a;
        endcase
    end else begin
        sbox_kout_aes_256_clk_a = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_a = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_a = 128'h0;
        case (clk_cnt_all)
            6'ha: begin
                sbox_dout_aes_256_clk_a[127:120] = AES_256_out_4;
                sbox_dout_aes_256_clk_a[119:112] = AES_256_out_5;
                sbox_dout_aes_256_clk_a[111:104] = AES_256_out_6;
                sbox_dout_aes_256_clk_a[103:96]  = AES_256_out_7;
                sbox_dout_aes_256_clk_a[95:88]   = AES_256_out_8;
                sbox_dout_aes_256_clk_a[87:80]   = AES_256_out_9;
                sbox_dout_aes_256_clk_a[79:72]   = AES_256_out_10;
                sbox_dout_aes_256_clk_a[71:64]   = AES_256_out_11;
                sbox_dout_aes_256_clk_a[63:56]   = AES_256_out_12;
                sbox_dout_aes_256_clk_a[55:48]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_a = sbox_dout_aes_256_clk_a;
        endcase
    end else begin
        sbox_dout_aes_256_clk_a = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_b = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_b = 128'h0;
        case (clk_cnt_all)
            6'hb: begin
                sbox_dout_aes_256_clk_b[47:40]   = AES_256_out_0;
                sbox_dout_aes_256_clk_b[39:32]   = AES_256_out_1;
                sbox_dout_aes_256_clk_b[31:24]   = AES_256_out_2;
                sbox_dout_aes_256_clk_b[23:16]   = AES_256_out_3;
                sbox_dout_aes_256_clk_b[15:8]    = AES_256_out_4;
                sbox_dout_aes_256_clk_b[7:0]     = AES_256_out_5;
                sbox_dout_aes_256_clk_b[127:120] = AES_256_out_10;
                sbox_dout_aes_256_clk_b[119:112] = AES_256_out_11;
                sbox_dout_aes_256_clk_b[111:104] = AES_256_out_12;
                sbox_dout_aes_256_clk_b[103:96]  = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_b = sbox_dout_aes_256_clk_b;
        endcase
    end else begin
        sbox_dout_aes_256_clk_b = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_b = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_b = 32'h0;
        case (clk_cnt_all)
            6'hb: begin
                sbox_kout_aes_256_clk_b[31:24]   = AES_256_out_6;
                sbox_kout_aes_256_clk_b[23:16]   = AES_256_out_7;
                sbox_kout_aes_256_clk_b[15:8]    = AES_256_out_8;
                sbox_kout_aes_256_clk_b[7:0]     = AES_256_out_9;
            end
            default: sbox_kout_aes_256_clk_b = sbox_kout_aes_256_clk_b;
        endcase
    end else begin
        sbox_kout_aes_256_clk_b = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_c = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_c = 128'h0;
        case (clk_cnt_all)
            6'hc: begin
                sbox_dout_aes_256_clk_c[95:88]   = AES_256_out_0;
                sbox_dout_aes_256_clk_c[87:80]   = AES_256_out_1;
                sbox_dout_aes_256_clk_c[79:72]   = AES_256_out_2;
                sbox_dout_aes_256_clk_c[71:64]   = AES_256_out_3;
                sbox_dout_aes_256_clk_c[63:56]   = AES_256_out_4;
                sbox_dout_aes_256_clk_c[55:48]   = AES_256_out_5;
                sbox_dout_aes_256_clk_c[47:40]   = AES_256_out_6;
                sbox_dout_aes_256_clk_c[39:32]   = AES_256_out_7;
                sbox_dout_aes_256_clk_c[31:24]   = AES_256_out_8;
                sbox_dout_aes_256_clk_c[23:16]   = AES_256_out_9;
                sbox_dout_aes_256_clk_c[15:8]    = AES_256_out_10;
                sbox_dout_aes_256_clk_c[7:0]     = AES_256_out_11;
            end
            default: sbox_dout_aes_256_clk_c = sbox_dout_aes_256_clk_c;
        endcase
    end else begin
        sbox_dout_aes_256_clk_c = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_c = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_c = 32'h0;
        case (clk_cnt_all)
            6'hc: begin
                sbox_kout_aes_256_clk_c[31:24]   = AES_256_out_12;
                sbox_kout_aes_256_clk_c[23:16]   = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_c = sbox_kout_aes_256_clk_c;
        endcase
    end else begin
        sbox_kout_aes_256_clk_c = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_d = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_d = 32'h0;
        case (clk_cnt_all)
            6'hd: begin
                sbox_kout_aes_256_clk_d[15:8]    = AES_256_out_0;
                sbox_kout_aes_256_clk_d[7:0]     = AES_256_out_1;
            end
            default: sbox_kout_aes_256_clk_d = sbox_kout_aes_256_clk_d;
        endcase
    end else begin
        sbox_kout_aes_256_clk_d = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_d = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_d = 128'h0;
        case (clk_cnt_all)
            6'hd: begin
                sbox_dout_aes_256_clk_d[127:120] = AES_256_out_2;
                sbox_dout_aes_256_clk_d[119:112] = AES_256_out_3;
                sbox_dout_aes_256_clk_d[111:104] = AES_256_out_4;
                sbox_dout_aes_256_clk_d[103:96]  = AES_256_out_5;
                sbox_dout_aes_256_clk_d[95:88]   = AES_256_out_6;
                sbox_dout_aes_256_clk_d[87:80]   = AES_256_out_7;
                sbox_dout_aes_256_clk_d[79:72]   = AES_256_out_8;
                sbox_dout_aes_256_clk_d[71:64]   = AES_256_out_9;
                sbox_dout_aes_256_clk_d[63:56]   = AES_256_out_10;
                sbox_dout_aes_256_clk_d[55:48]   = AES_256_out_11;
                sbox_dout_aes_256_clk_d[47:40]   = AES_256_out_12;
                sbox_dout_aes_256_clk_d[39:32]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_d = sbox_dout_aes_256_clk_d;
        endcase
    end else begin
        sbox_dout_aes_256_clk_d = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_e = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_e = 128'h0;
        case (clk_cnt_all)
            6'he: begin
                sbox_dout_aes_256_clk_e[31:24]   = AES_256_out_0;
                sbox_dout_aes_256_clk_e[23:16]   = AES_256_out_1;
                sbox_dout_aes_256_clk_e[15:8]    = AES_256_out_2;
                sbox_dout_aes_256_clk_e[7:0]     = AES_256_out_3;
                sbox_dout_aes_256_clk_e[127:120] = AES_256_out_8;
                sbox_dout_aes_256_clk_e[119:112] = AES_256_out_9;
                sbox_dout_aes_256_clk_e[111:104] = AES_256_out_10;
                sbox_dout_aes_256_clk_e[103:96]  = AES_256_out_11;
                sbox_dout_aes_256_clk_e[95:88]   = AES_256_out_12;
                sbox_dout_aes_256_clk_e[87:80]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_e = sbox_dout_aes_256_clk_e;
        endcase
    end else begin
        sbox_dout_aes_256_clk_e = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_e = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_e = 32'h0;
        case (clk_cnt_all)
            6'he: begin
                sbox_kout_aes_256_clk_e[31:24]   = AES_256_out_4;
                sbox_kout_aes_256_clk_e[23:16]   = AES_256_out_5;
                sbox_kout_aes_256_clk_e[15:8]    = AES_256_out_6;
                sbox_kout_aes_256_clk_e[7:0]     = AES_256_out_7;
            end
            default: sbox_kout_aes_256_clk_e = sbox_kout_aes_256_clk_e;
        endcase
    end else begin
        sbox_kout_aes_256_clk_e = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_f = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_f = 128'h0;
        case (clk_cnt_all)
            6'hf: begin
                sbox_dout_aes_256_clk_f[79:72]   = AES_256_out_0;
                sbox_dout_aes_256_clk_f[71:64]   = AES_256_out_1;
                sbox_dout_aes_256_clk_f[63:56]   = AES_256_out_2;
                sbox_dout_aes_256_clk_f[55:48]   = AES_256_out_3;
                sbox_dout_aes_256_clk_f[47:40]   = AES_256_out_4;
                sbox_dout_aes_256_clk_f[39:32]   = AES_256_out_5;
                sbox_dout_aes_256_clk_f[31:24]   = AES_256_out_6;
                sbox_dout_aes_256_clk_f[23:16]   = AES_256_out_7;
                sbox_dout_aes_256_clk_f[15:8]    = AES_256_out_8;
                sbox_dout_aes_256_clk_f[7:0]     = AES_256_out_9;
            end
            default: sbox_dout_aes_256_clk_f = sbox_dout_aes_256_clk_f;
        endcase
    end else begin
        sbox_dout_aes_256_clk_f = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_f = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_f = 32'h0;
        case (clk_cnt_all)
            6'hf: begin
                sbox_kout_aes_256_clk_f[31:24]   = AES_256_out_10;
                sbox_kout_aes_256_clk_f[23:16]   = AES_256_out_11;
                sbox_kout_aes_256_clk_f[15:8]    = AES_256_out_12;
                sbox_kout_aes_256_clk_f[7:0]     = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_f = sbox_kout_aes_256_clk_f;
        endcase
    end else begin
        sbox_kout_aes_256_clk_f = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_10 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_10 = 128'h0;
        case (clk_cnt_all)
            6'h10: begin
                sbox_dout_aes_256_clk_10[127:120] = AES_256_out_0;
                sbox_dout_aes_256_clk_10[119:112] = AES_256_out_1;
                sbox_dout_aes_256_clk_10[111:104] = AES_256_out_2;
                sbox_dout_aes_256_clk_10[103:96]  = AES_256_out_3;
                sbox_dout_aes_256_clk_10[95:88]   = AES_256_out_4;
                sbox_dout_aes_256_clk_10[87:80]   = AES_256_out_5;
                sbox_dout_aes_256_clk_10[79:72]   = AES_256_out_6;
                sbox_dout_aes_256_clk_10[71:64]   = AES_256_out_7;
                sbox_dout_aes_256_clk_10[63:56]   = AES_256_out_8;
                sbox_dout_aes_256_clk_10[55:48]   = AES_256_out_9;
                sbox_dout_aes_256_clk_10[47:40]   = AES_256_out_10;
                sbox_dout_aes_256_clk_10[39:32]   = AES_256_out_11;
                sbox_dout_aes_256_clk_10[31:24]   = AES_256_out_12;
                sbox_dout_aes_256_clk_10[23:16]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_10 = sbox_dout_aes_256_clk_10;
        endcase
    end else begin
        sbox_dout_aes_256_clk_10 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_11 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_11 = 128'h0;
        case (clk_cnt_all)
            6'h11: begin
                sbox_dout_aes_256_clk_11[15:8]    = AES_256_out_0;
                sbox_dout_aes_256_clk_11[7:0]     = AES_256_out_1;
                sbox_dout_aes_256_clk_11[127:120] = AES_256_out_6;
                sbox_dout_aes_256_clk_11[119:112] = AES_256_out_7;
                sbox_dout_aes_256_clk_11[111:104] = AES_256_out_8;
                sbox_dout_aes_256_clk_11[103:96]  = AES_256_out_9;
                sbox_dout_aes_256_clk_11[95:88]   = AES_256_out_10;
                sbox_dout_aes_256_clk_11[87:80]   = AES_256_out_11;
                sbox_dout_aes_256_clk_11[79:72]   = AES_256_out_12;
                sbox_dout_aes_256_clk_11[71:64]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_11 = sbox_dout_aes_256_clk_11;
        endcase
    end else begin
        sbox_dout_aes_256_clk_11 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_11 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_11 = 32'h0;
        case (clk_cnt_all)
            6'h11: begin
                sbox_kout_aes_256_clk_11[31:24]   = AES_256_out_2;
                sbox_kout_aes_256_clk_11[23:16]   = AES_256_out_3;
                sbox_kout_aes_256_clk_11[15:8]    = AES_256_out_4;
                sbox_kout_aes_256_clk_11[7:0]     = AES_256_out_5;
            end
            default: sbox_kout_aes_256_clk_11 = sbox_kout_aes_256_clk_11;
        endcase
    end else begin
        sbox_kout_aes_256_clk_11 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_12 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_12 = 128'h0;
        case (clk_cnt_all)
            6'h12: begin
                sbox_dout_aes_256_clk_12[63:56]   = AES_256_out_0;
                sbox_dout_aes_256_clk_12[55:48]   = AES_256_out_1;
                sbox_dout_aes_256_clk_12[47:40]   = AES_256_out_2;
                sbox_dout_aes_256_clk_12[39:32]   = AES_256_out_3;
                sbox_dout_aes_256_clk_12[31:24]   = AES_256_out_4;
                sbox_dout_aes_256_clk_12[23:16]   = AES_256_out_5;
                sbox_dout_aes_256_clk_12[15:8]    = AES_256_out_6;
                sbox_dout_aes_256_clk_12[7:0]     = AES_256_out_7;
                sbox_dout_aes_256_clk_12[127:120] = AES_256_out_12;
                sbox_dout_aes_256_clk_12[119:112] = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_12 = sbox_dout_aes_256_clk_12;
        endcase
    end else begin
        sbox_dout_aes_256_clk_12 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_12 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_12 = 32'h0;
        case (clk_cnt_all)
            6'h12: begin
                sbox_kout_aes_256_clk_12[31:24]   = AES_256_out_8;
                sbox_kout_aes_256_clk_12[23:16]   = AES_256_out_9;
                sbox_kout_aes_256_clk_12[15:8]    = AES_256_out_10;
                sbox_kout_aes_256_clk_12[7:0]     = AES_256_out_11;
            end
            default: sbox_kout_aes_256_clk_12 = sbox_kout_aes_256_clk_12;
        endcase
    end else begin
        sbox_kout_aes_256_clk_12 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_13 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_13 = 128'h0;
        case (clk_cnt_all)
            6'h13: begin
                sbox_dout_aes_256_clk_13[111:104] = AES_256_out_0;
                sbox_dout_aes_256_clk_13[103:96]  = AES_256_out_1;
                sbox_dout_aes_256_clk_13[95:88]   = AES_256_out_2;
                sbox_dout_aes_256_clk_13[87:80]   = AES_256_out_3;
                sbox_dout_aes_256_clk_13[79:72]   = AES_256_out_4;
                sbox_dout_aes_256_clk_13[71:64]   = AES_256_out_5;
                sbox_dout_aes_256_clk_13[63:56]   = AES_256_out_6;
                sbox_dout_aes_256_clk_13[55:48]   = AES_256_out_7;
                sbox_dout_aes_256_clk_13[47:40]   = AES_256_out_8;
                sbox_dout_aes_256_clk_13[39:32]   = AES_256_out_9;
                sbox_dout_aes_256_clk_13[31:24]   = AES_256_out_10;
                sbox_dout_aes_256_clk_13[23:16]   = AES_256_out_11;
                sbox_dout_aes_256_clk_13[15:8]    = AES_256_out_12;
                sbox_dout_aes_256_clk_13[7:0]     = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_13 = sbox_dout_aes_256_clk_13;
        endcase
    end else begin
        sbox_dout_aes_256_clk_13 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_14 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_14 = 32'h0;
        case (clk_cnt_all)
            6'h14: begin
                sbox_kout_aes_256_clk_14[31:24]   = AES_256_out_0;
                sbox_kout_aes_256_clk_14[23:16]   = AES_256_out_1;
                sbox_kout_aes_256_clk_14[15:8 ]   = AES_256_out_2;
                sbox_kout_aes_256_clk_14[7:0]     = AES_256_out_3;
            end
            default: sbox_kout_aes_256_clk_14 = sbox_kout_aes_256_clk_14;
        endcase
    end else begin
        sbox_kout_aes_256_clk_14 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_14 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_14 = 128'h0;
        case (clk_cnt_all)
            6'h14: begin
                sbox_dout_aes_256_clk_14[127:120] = AES_256_out_4;
                sbox_dout_aes_256_clk_14[119:112] = AES_256_out_5;
                sbox_dout_aes_256_clk_14[111:104] = AES_256_out_6;
                sbox_dout_aes_256_clk_14[103:96]  = AES_256_out_7;
                sbox_dout_aes_256_clk_14[95:88]   = AES_256_out_8;
                sbox_dout_aes_256_clk_14[87:80]   = AES_256_out_9;
                sbox_dout_aes_256_clk_14[79:72]   = AES_256_out_10;
                sbox_dout_aes_256_clk_14[71:64]   = AES_256_out_11;
                sbox_dout_aes_256_clk_14[63:56]   = AES_256_out_12;
                sbox_dout_aes_256_clk_14[55:48]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_14 = sbox_dout_aes_256_clk_14;
        endcase
    end else begin
        sbox_dout_aes_256_clk_14 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_15 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_15 = 128'h0;
        case (clk_cnt_all)
            6'h15: begin
                sbox_dout_aes_256_clk_15[47:40]   = AES_256_out_0;
                sbox_dout_aes_256_clk_15[39:32]   = AES_256_out_1;
                sbox_dout_aes_256_clk_15[31:24]   = AES_256_out_2;
                sbox_dout_aes_256_clk_15[23:16]   = AES_256_out_3;
                sbox_dout_aes_256_clk_15[15:8]    = AES_256_out_4;
                sbox_dout_aes_256_clk_15[7:0]     = AES_256_out_5;
                sbox_dout_aes_256_clk_15[127:120] = AES_256_out_10;
                sbox_dout_aes_256_clk_15[119:112] = AES_256_out_11;
                sbox_dout_aes_256_clk_15[111:104] = AES_256_out_12;
                sbox_dout_aes_256_clk_15[103:96]  = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_15 = sbox_dout_aes_256_clk_15;
        endcase
    end else begin
        sbox_dout_aes_256_clk_15 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_15 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_15 = 32'h0;
        case (clk_cnt_all)
            6'h15: begin
                sbox_kout_aes_256_clk_15[31:24]   = AES_256_out_6;
                sbox_kout_aes_256_clk_15[23:16]   = AES_256_out_7;
                sbox_kout_aes_256_clk_15[15:8]    = AES_256_out_8;
                sbox_kout_aes_256_clk_15[7:0]     = AES_256_out_9;
            end
            default: sbox_kout_aes_256_clk_15 = sbox_kout_aes_256_clk_15;
        endcase
    end else begin
        sbox_kout_aes_256_clk_15 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_16 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_16 = 128'h0;
        case (clk_cnt_all)
            6'h16: begin
                sbox_dout_aes_256_clk_16[95:88]   = AES_256_out_0;
                sbox_dout_aes_256_clk_16[87:80]   = AES_256_out_1;
                sbox_dout_aes_256_clk_16[79:72]   = AES_256_out_2;
                sbox_dout_aes_256_clk_16[71:64]   = AES_256_out_3;
                sbox_dout_aes_256_clk_16[63:56]   = AES_256_out_4;
                sbox_dout_aes_256_clk_16[55:48]   = AES_256_out_5;
                sbox_dout_aes_256_clk_16[47:40]   = AES_256_out_6;
                sbox_dout_aes_256_clk_16[39:32]   = AES_256_out_7;
                sbox_dout_aes_256_clk_16[31:24]   = AES_256_out_8;
                sbox_dout_aes_256_clk_16[23:16]   = AES_256_out_9;
                sbox_dout_aes_256_clk_16[15:8]    = AES_256_out_10;
                sbox_dout_aes_256_clk_16[7:0]     = AES_256_out_11;
            end
            default: sbox_dout_aes_256_clk_16 = sbox_dout_aes_256_clk_16;
        endcase
    end else begin
        sbox_dout_aes_256_clk_16 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_16 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_16 = 32'h0;
        case (clk_cnt_all)
            6'h16: begin
                sbox_kout_aes_256_clk_16[31:24]   = AES_256_out_12;
                sbox_kout_aes_256_clk_16[23:16]   = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_16 = sbox_kout_aes_256_clk_16;
        endcase
    end else begin
        sbox_kout_aes_256_clk_16 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_17 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_17 = 32'h0;
        case (clk_cnt_all)
            6'h17: begin
                sbox_kout_aes_256_clk_17[15:8]    = AES_256_out_0;
                sbox_kout_aes_256_clk_17[7:0]     = AES_256_out_1;
            end
            default: sbox_kout_aes_256_clk_17 = sbox_kout_aes_256_clk_17;
        endcase
    end else begin
        sbox_kout_aes_256_clk_17 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_17 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_17 = 128'h0;
        case (clk_cnt_all)
            6'h17: begin
                sbox_dout_aes_256_clk_17[127:120] = AES_256_out_2;
                sbox_dout_aes_256_clk_17[119:112] = AES_256_out_3;
                sbox_dout_aes_256_clk_17[111:104] = AES_256_out_4;
                sbox_dout_aes_256_clk_17[103:96]  = AES_256_out_5;
                sbox_dout_aes_256_clk_17[95:88]   = AES_256_out_6;
                sbox_dout_aes_256_clk_17[87:80]   = AES_256_out_7;
                sbox_dout_aes_256_clk_17[79:72]   = AES_256_out_8;
                sbox_dout_aes_256_clk_17[71:64]   = AES_256_out_9;
                sbox_dout_aes_256_clk_17[63:56]   = AES_256_out_10;
                sbox_dout_aes_256_clk_17[55:48]   = AES_256_out_11;
                sbox_dout_aes_256_clk_17[47:40]   = AES_256_out_12;
                sbox_dout_aes_256_clk_17[39:32]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_17 = sbox_dout_aes_256_clk_17;
        endcase
    end else begin
        sbox_dout_aes_256_clk_17 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_18 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_18 = 128'h0;
        case (clk_cnt_all)
            6'h18: begin
                sbox_dout_aes_256_clk_18[31:24]   = AES_256_out_0;
                sbox_dout_aes_256_clk_18[23:16]   = AES_256_out_1;
                sbox_dout_aes_256_clk_18[15:8]    = AES_256_out_2;
                sbox_dout_aes_256_clk_18[7:0]     = AES_256_out_3;
                sbox_dout_aes_256_clk_18[127:120] = AES_256_out_8;
                sbox_dout_aes_256_clk_18[119:112] = AES_256_out_9;
                sbox_dout_aes_256_clk_18[111:104] = AES_256_out_10;
                sbox_dout_aes_256_clk_18[103:96]  = AES_256_out_11;
                sbox_dout_aes_256_clk_18[95:88]   = AES_256_out_12;
                sbox_dout_aes_256_clk_18[87:80]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_18 = sbox_dout_aes_256_clk_18;
        endcase
    end else begin
        sbox_dout_aes_256_clk_18 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_18 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_18 = 32'h0;
        case (clk_cnt_all)
            6'h18: begin
                sbox_kout_aes_256_clk_18[31:24]   = AES_256_out_4;
                sbox_kout_aes_256_clk_18[23:16]   = AES_256_out_5;
                sbox_kout_aes_256_clk_18[15:8]    = AES_256_out_6;
                sbox_kout_aes_256_clk_18[7:0]     = AES_256_out_7;
            end
            default: sbox_kout_aes_256_clk_18 = sbox_kout_aes_256_clk_18;
        endcase
    end else begin
        sbox_kout_aes_256_clk_18 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_19 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_19 = 128'h0;
        case (clk_cnt_all)
            6'h19: begin
                sbox_dout_aes_256_clk_19[79:72]   = AES_256_out_0;
                sbox_dout_aes_256_clk_19[71:64]   = AES_256_out_1;
                sbox_dout_aes_256_clk_19[63:56]   = AES_256_out_2;
                sbox_dout_aes_256_clk_19[55:48]   = AES_256_out_3;
                sbox_dout_aes_256_clk_19[47:40]   = AES_256_out_4;
                sbox_dout_aes_256_clk_19[39:32]   = AES_256_out_5;
                sbox_dout_aes_256_clk_19[31:24]   = AES_256_out_6;
                sbox_dout_aes_256_clk_19[23:16]   = AES_256_out_7;
                sbox_dout_aes_256_clk_19[15:8]    = AES_256_out_8;
                sbox_dout_aes_256_clk_19[7:0]     = AES_256_out_9;
            end
            default: sbox_dout_aes_256_clk_19 = sbox_dout_aes_256_clk_19;
        endcase
    end else begin
        sbox_dout_aes_256_clk_19 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_19 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_19 = 32'h0;
        case (clk_cnt_all)
            6'h19: begin
                sbox_kout_aes_256_clk_19[31:24]   = AES_256_out_10;
                sbox_kout_aes_256_clk_19[23:16]   = AES_256_out_11;
                sbox_kout_aes_256_clk_19[15:8]    = AES_256_out_12;
                sbox_kout_aes_256_clk_19[7:0]     = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_19 = sbox_kout_aes_256_clk_19;
        endcase
    end else begin
        sbox_kout_aes_256_clk_19 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_1a = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_1a = 128'h0;
        case (clk_cnt_all)
            6'h1a: begin
                sbox_dout_aes_256_clk_1a[127:120] = AES_256_out_0;
                sbox_dout_aes_256_clk_1a[119:112] = AES_256_out_1;
                sbox_dout_aes_256_clk_1a[111:104] = AES_256_out_2;
                sbox_dout_aes_256_clk_1a[103:96]  = AES_256_out_3;
                sbox_dout_aes_256_clk_1a[95:88]   = AES_256_out_4;
                sbox_dout_aes_256_clk_1a[87:80]   = AES_256_out_5;
                sbox_dout_aes_256_clk_1a[79:72]   = AES_256_out_6;
                sbox_dout_aes_256_clk_1a[71:64]   = AES_256_out_7;
                sbox_dout_aes_256_clk_1a[63:56]   = AES_256_out_8;
                sbox_dout_aes_256_clk_1a[55:48]   = AES_256_out_9;
                sbox_dout_aes_256_clk_1a[47:40]   = AES_256_out_10;
                sbox_dout_aes_256_clk_1a[39:32]   = AES_256_out_11;
                sbox_dout_aes_256_clk_1a[31:24]   = AES_256_out_12;
                sbox_dout_aes_256_clk_1a[23:16]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_1a = sbox_dout_aes_256_clk_1a;
        endcase
    end else begin
        sbox_dout_aes_256_clk_1a = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_1b = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_1b = 128'h0;
        case (clk_cnt_all)
            6'h1b: begin
                sbox_dout_aes_256_clk_1b[15:8]    = AES_256_out_0;
                sbox_dout_aes_256_clk_1b[7:0]     = AES_256_out_1;
                sbox_dout_aes_256_clk_1b[127:120] = AES_256_out_6;
                sbox_dout_aes_256_clk_1b[119:112] = AES_256_out_7;
                sbox_dout_aes_256_clk_1b[111:104] = AES_256_out_8;
                sbox_dout_aes_256_clk_1b[103:96]  = AES_256_out_9;
                sbox_dout_aes_256_clk_1b[95:88]   = AES_256_out_10;
                sbox_dout_aes_256_clk_1b[87:80]   = AES_256_out_11;
                sbox_dout_aes_256_clk_1b[79:72]   = AES_256_out_12;
                sbox_dout_aes_256_clk_1b[71:64]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_1b = sbox_dout_aes_256_clk_1b;
        endcase
    end else begin
        sbox_dout_aes_256_clk_1b = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_1b = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_1b = 32'h0;
        case (clk_cnt_all)
            6'h1b: begin
                sbox_kout_aes_256_clk_1b[31:24]   = AES_256_out_2;
                sbox_kout_aes_256_clk_1b[23:16]   = AES_256_out_3;
                sbox_kout_aes_256_clk_1b[15:8]    = AES_256_out_4;
                sbox_kout_aes_256_clk_1b[7:0]     = AES_256_out_5;
            end
            default: sbox_kout_aes_256_clk_1b = sbox_kout_aes_256_clk_1b;
        endcase
    end else begin
        sbox_kout_aes_256_clk_1b = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_1c = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_1c = 128'h0;
        case (clk_cnt_all)
            6'h1c: begin
                sbox_dout_aes_256_clk_1c[63:56]   = AES_256_out_0;
                sbox_dout_aes_256_clk_1c[55:48]   = AES_256_out_1;
                sbox_dout_aes_256_clk_1c[47:40]   = AES_256_out_2;
                sbox_dout_aes_256_clk_1c[39:32]   = AES_256_out_3;
                sbox_dout_aes_256_clk_1c[31:24]   = AES_256_out_4;
                sbox_dout_aes_256_clk_1c[23:16]   = AES_256_out_5;
                sbox_dout_aes_256_clk_1c[15:8]    = AES_256_out_6;
                sbox_dout_aes_256_clk_1c[7:0]     = AES_256_out_7;
                sbox_dout_aes_256_clk_1c[127:120] = AES_256_out_12;
                sbox_dout_aes_256_clk_1c[119:112] = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_1c = sbox_dout_aes_256_clk_1c;
        endcase
    end else begin
        sbox_dout_aes_256_clk_1c = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_1c = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_1c = 32'h0;
        case (clk_cnt_all)
            6'h1c: begin
                sbox_kout_aes_256_clk_1c[31:24]   = AES_256_out_8;
                sbox_kout_aes_256_clk_1c[23:16]   = AES_256_out_9;
                sbox_kout_aes_256_clk_1c[15:8]    = AES_256_out_10;
                sbox_kout_aes_256_clk_1c[7:0]     = AES_256_out_11;
            end
            default: sbox_kout_aes_256_clk_1c = sbox_kout_aes_256_clk_1c;
        endcase
    end else begin
        sbox_kout_aes_256_clk_1c = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_1d = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_1d = 128'h0;
        case (clk_cnt_all)
            6'h1d: begin
                sbox_dout_aes_256_clk_1d[111:104] = AES_256_out_0;
                sbox_dout_aes_256_clk_1d[103:96]  = AES_256_out_1;
                sbox_dout_aes_256_clk_1d[95:88]   = AES_256_out_2;
                sbox_dout_aes_256_clk_1d[87:80]   = AES_256_out_3;
                sbox_dout_aes_256_clk_1d[79:72]   = AES_256_out_4;
                sbox_dout_aes_256_clk_1d[71:64]   = AES_256_out_5;
                sbox_dout_aes_256_clk_1d[63:56]   = AES_256_out_6;
                sbox_dout_aes_256_clk_1d[55:48]   = AES_256_out_7;
                sbox_dout_aes_256_clk_1d[47:40]   = AES_256_out_8;
                sbox_dout_aes_256_clk_1d[39:32]   = AES_256_out_9;
                sbox_dout_aes_256_clk_1d[31:24]   = AES_256_out_10;
                sbox_dout_aes_256_clk_1d[23:16]   = AES_256_out_11;
                sbox_dout_aes_256_clk_1d[15:8]    = AES_256_out_12;
                sbox_dout_aes_256_clk_1d[7:0]     = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_1d = sbox_dout_aes_256_clk_1d;
        endcase
    end else begin
        sbox_dout_aes_256_clk_1d = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_1e = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_1e = 32'h0;
        case (clk_cnt_all)
            6'h1e: begin
                sbox_kout_aes_256_clk_1e[31:24]   = AES_256_out_0;
                sbox_kout_aes_256_clk_1e[23:16]   = AES_256_out_1;
                sbox_kout_aes_256_clk_1e[15:8 ]   = AES_256_out_2;
                sbox_kout_aes_256_clk_1e[7:0]     = AES_256_out_3;
            end
            default: sbox_kout_aes_256_clk_1e = sbox_kout_aes_256_clk_1e;
        endcase
    end else begin
        sbox_kout_aes_256_clk_1e = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_1e = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_1e = 128'h0;
        case (clk_cnt_all)
            6'h1e: begin
                sbox_dout_aes_256_clk_1e[127:120] = AES_256_out_4;
                sbox_dout_aes_256_clk_1e[119:112] = AES_256_out_5;
                sbox_dout_aes_256_clk_1e[111:104] = AES_256_out_6;
                sbox_dout_aes_256_clk_1e[103:96]  = AES_256_out_7;
                sbox_dout_aes_256_clk_1e[95:88]   = AES_256_out_8;
                sbox_dout_aes_256_clk_1e[87:80]   = AES_256_out_9;
                sbox_dout_aes_256_clk_1e[79:72]   = AES_256_out_10;
                sbox_dout_aes_256_clk_1e[71:64]   = AES_256_out_11;
                sbox_dout_aes_256_clk_1e[63:56]   = AES_256_out_12;
                sbox_dout_aes_256_clk_1e[55:48]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_1e = sbox_dout_aes_256_clk_1e;
        endcase
    end else begin
        sbox_dout_aes_256_clk_1e = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_1f = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_1f = 128'h0;
        case (clk_cnt_all)
            6'h1f: begin
                sbox_dout_aes_256_clk_1f[47:40]   = AES_256_out_0;
                sbox_dout_aes_256_clk_1f[39:32]   = AES_256_out_1;
                sbox_dout_aes_256_clk_1f[31:24]   = AES_256_out_2;
                sbox_dout_aes_256_clk_1f[23:16]   = AES_256_out_3;
                sbox_dout_aes_256_clk_1f[15:8]    = AES_256_out_4;
                sbox_dout_aes_256_clk_1f[7:0]     = AES_256_out_5;
                sbox_dout_aes_256_clk_1f[127:120] = AES_256_out_10;
                sbox_dout_aes_256_clk_1f[119:112] = AES_256_out_11;
                sbox_dout_aes_256_clk_1f[111:104] = AES_256_out_12;
                sbox_dout_aes_256_clk_1f[103:96]  = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_1f = sbox_dout_aes_256_clk_1f;
        endcase
    end else begin
        sbox_dout_aes_256_clk_1f = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_1f = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_1f = 32'h0;
        case (clk_cnt_all)
            6'h1f: begin
                sbox_kout_aes_256_clk_1f[31:24]   = AES_256_out_6;
                sbox_kout_aes_256_clk_1f[23:16]   = AES_256_out_7;
                sbox_kout_aes_256_clk_1f[15:8]    = AES_256_out_8;
                sbox_kout_aes_256_clk_1f[7:0]     = AES_256_out_9;
            end
            default: sbox_kout_aes_256_clk_1f = sbox_kout_aes_256_clk_1f;
        endcase
    end else begin
        sbox_kout_aes_256_clk_1f = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_20 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_20 = 128'h0;
        case (clk_cnt_all)
            6'h20: begin
                sbox_dout_aes_256_clk_20[95:88]   = AES_256_out_0;
                sbox_dout_aes_256_clk_20[87:80]   = AES_256_out_1;
                sbox_dout_aes_256_clk_20[79:72]   = AES_256_out_2;
                sbox_dout_aes_256_clk_20[71:64]   = AES_256_out_3;
                sbox_dout_aes_256_clk_20[63:56]   = AES_256_out_4;
                sbox_dout_aes_256_clk_20[55:48]   = AES_256_out_5;
                sbox_dout_aes_256_clk_20[47:40]   = AES_256_out_6;
                sbox_dout_aes_256_clk_20[39:32]   = AES_256_out_7;
                sbox_dout_aes_256_clk_20[31:24]   = AES_256_out_8;
                sbox_dout_aes_256_clk_20[23:16]   = AES_256_out_9;
                sbox_dout_aes_256_clk_20[15:8]    = AES_256_out_10;
                sbox_dout_aes_256_clk_20[7:0]     = AES_256_out_11;
            end
            default: sbox_dout_aes_256_clk_20 = sbox_dout_aes_256_clk_20;
        endcase
    end else begin
        sbox_dout_aes_256_clk_20 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_20 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_20 = 32'h0;
        case (clk_cnt_all)
            6'h20: begin
                sbox_kout_aes_256_clk_20[31:24]   = AES_256_out_12;
                sbox_kout_aes_256_clk_20[23:16]   = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_20 = sbox_kout_aes_256_clk_20;
        endcase
    end else begin
        sbox_kout_aes_256_clk_20 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_21 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_21 = 32'h0;
        case (clk_cnt_all)
            6'h21: begin
                sbox_kout_aes_256_clk_21[15:8]    = AES_256_out_0;
                sbox_kout_aes_256_clk_21[7:0]     = AES_256_out_1;
            end
            default: sbox_kout_aes_256_clk_21 = sbox_kout_aes_256_clk_21;
        endcase
    end else begin
        sbox_kout_aes_256_clk_21 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_21 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_21 = 128'h0;
        case (clk_cnt_all)
            6'h21: begin
                sbox_dout_aes_256_clk_21[127:120] = AES_256_out_2;
                sbox_dout_aes_256_clk_21[119:112] = AES_256_out_3;
                sbox_dout_aes_256_clk_21[111:104] = AES_256_out_4;
                sbox_dout_aes_256_clk_21[103:96]  = AES_256_out_5;
                sbox_dout_aes_256_clk_21[95:88]   = AES_256_out_6;
                sbox_dout_aes_256_clk_21[87:80]   = AES_256_out_7;
                sbox_dout_aes_256_clk_21[79:72]   = AES_256_out_8;
                sbox_dout_aes_256_clk_21[71:64]   = AES_256_out_9;
                sbox_dout_aes_256_clk_21[63:56]   = AES_256_out_10;
                sbox_dout_aes_256_clk_21[55:48]   = AES_256_out_11;
                sbox_dout_aes_256_clk_21[47:40]   = AES_256_out_12;
                sbox_dout_aes_256_clk_21[39:32]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_21 = sbox_dout_aes_256_clk_21;
        endcase
    end else begin
        sbox_dout_aes_256_clk_21 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_22 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_22 = 128'h0;
        case (clk_cnt_all)
            6'h22: begin
                sbox_dout_aes_256_clk_22[31:24]   = AES_256_out_0;
                sbox_dout_aes_256_clk_22[23:16]   = AES_256_out_1;
                sbox_dout_aes_256_clk_22[15:8]    = AES_256_out_2;
                sbox_dout_aes_256_clk_22[7:0]     = AES_256_out_3;
                sbox_dout_aes_256_clk_22[127:120] = AES_256_out_8;
                sbox_dout_aes_256_clk_22[119:112] = AES_256_out_9;
                sbox_dout_aes_256_clk_22[111:104] = AES_256_out_10;
                sbox_dout_aes_256_clk_22[103:96]  = AES_256_out_11;
                sbox_dout_aes_256_clk_22[95:88]   = AES_256_out_12;
                sbox_dout_aes_256_clk_22[87:80]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_22 = sbox_dout_aes_256_clk_22;
        endcase
    end else begin
        sbox_dout_aes_256_clk_22 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_22 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_22 = 32'h0;
        case (clk_cnt_all)
            6'h22: begin
                sbox_kout_aes_256_clk_22[31:24]   = AES_256_out_4;
                sbox_kout_aes_256_clk_22[23:16]   = AES_256_out_5;
                sbox_kout_aes_256_clk_22[15:8]    = AES_256_out_6;
                sbox_kout_aes_256_clk_22[7:0]     = AES_256_out_7;
            end
            default: sbox_kout_aes_256_clk_22 = sbox_kout_aes_256_clk_22;
        endcase
    end else begin
        sbox_kout_aes_256_clk_22 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_23 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_23 = 128'h0;
        case (clk_cnt_all)
            6'h23: begin
                sbox_dout_aes_256_clk_23[79:72]   = AES_256_out_0;
                sbox_dout_aes_256_clk_23[71:64]   = AES_256_out_1;
                sbox_dout_aes_256_clk_23[63:56]   = AES_256_out_2;
                sbox_dout_aes_256_clk_23[55:48]   = AES_256_out_3;
                sbox_dout_aes_256_clk_23[47:40]   = AES_256_out_4;
                sbox_dout_aes_256_clk_23[39:32]   = AES_256_out_5;
                sbox_dout_aes_256_clk_23[31:24]   = AES_256_out_6;
                sbox_dout_aes_256_clk_23[23:16]   = AES_256_out_7;
                sbox_dout_aes_256_clk_23[15:8]    = AES_256_out_8;
                sbox_dout_aes_256_clk_23[7:0]     = AES_256_out_9;
            end
            default: sbox_dout_aes_256_clk_23 = sbox_dout_aes_256_clk_23;
        endcase
    end else begin
        sbox_dout_aes_256_clk_23 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_23 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_23 = 32'h0;
        case (clk_cnt_all)
            6'h23: begin
                sbox_kout_aes_256_clk_23[31:24]   = AES_256_out_10;
                sbox_kout_aes_256_clk_23[23:16]   = AES_256_out_11;
                sbox_kout_aes_256_clk_23[15:8]    = AES_256_out_12;
                sbox_kout_aes_256_clk_23[7:0]     = AES_256_out_13;
            end
            default: sbox_kout_aes_256_clk_23 = sbox_kout_aes_256_clk_23;
        endcase
    end else begin
        sbox_kout_aes_256_clk_23 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_24 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_24 = 128'h0;
        case (clk_cnt_all)
            6'h24: begin
                sbox_dout_aes_256_clk_24[127:120] = AES_256_out_0;
                sbox_dout_aes_256_clk_24[119:112] = AES_256_out_1;
                sbox_dout_aes_256_clk_24[111:104] = AES_256_out_2;
                sbox_dout_aes_256_clk_24[103:96]  = AES_256_out_3;
                sbox_dout_aes_256_clk_24[95:88]   = AES_256_out_4;
                sbox_dout_aes_256_clk_24[87:80]   = AES_256_out_5;
                sbox_dout_aes_256_clk_24[79:72]   = AES_256_out_6;
                sbox_dout_aes_256_clk_24[71:64]   = AES_256_out_7;
                sbox_dout_aes_256_clk_24[63:56]   = AES_256_out_8;
                sbox_dout_aes_256_clk_24[55:48]   = AES_256_out_9;
                sbox_dout_aes_256_clk_24[47:40]   = AES_256_out_10;
                sbox_dout_aes_256_clk_24[39:32]   = AES_256_out_11;
                sbox_dout_aes_256_clk_24[31:24]   = AES_256_out_12;
                sbox_dout_aes_256_clk_24[23:16]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_24 = sbox_dout_aes_256_clk_24;
        endcase
    end else begin
        sbox_dout_aes_256_clk_24 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_25 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_25 = 128'h0;
        case (clk_cnt_all)
            6'h25: begin
                sbox_dout_aes_256_clk_25[15:8]    = AES_256_out_0;
                sbox_dout_aes_256_clk_25[7:0]     = AES_256_out_1;
                sbox_dout_aes_256_clk_25[127:120] = AES_256_out_6;
                sbox_dout_aes_256_clk_25[119:112] = AES_256_out_7;
                sbox_dout_aes_256_clk_25[111:104] = AES_256_out_8;
                sbox_dout_aes_256_clk_25[103:96]  = AES_256_out_9;
                sbox_dout_aes_256_clk_25[95:88]   = AES_256_out_10;
                sbox_dout_aes_256_clk_25[87:80]   = AES_256_out_11;
                sbox_dout_aes_256_clk_25[79:72]   = AES_256_out_12;
                sbox_dout_aes_256_clk_25[71:64]   = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_25 = sbox_dout_aes_256_clk_25;
        endcase
    end else begin
        sbox_dout_aes_256_clk_25 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_25 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_25 = 32'h0;
        case (clk_cnt_all)
            6'h25: begin
                sbox_kout_aes_256_clk_25[31:24]   = AES_256_out_2;
                sbox_kout_aes_256_clk_25[23:16]   = AES_256_out_3;
                sbox_kout_aes_256_clk_25[15:8]    = AES_256_out_4;
                sbox_kout_aes_256_clk_25[7:0]     = AES_256_out_5;
            end
            default: sbox_kout_aes_256_clk_25 = sbox_kout_aes_256_clk_25;
        endcase
    end else begin
        sbox_kout_aes_256_clk_25 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_26 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_26 = 128'h0;
        case (clk_cnt_all)
            6'h26: begin
                sbox_dout_aes_256_clk_26[63:56]   = AES_256_out_0;
                sbox_dout_aes_256_clk_26[55:48]   = AES_256_out_1;
                sbox_dout_aes_256_clk_26[47:40]   = AES_256_out_2;
                sbox_dout_aes_256_clk_26[39:32]   = AES_256_out_3;
                sbox_dout_aes_256_clk_26[31:24]   = AES_256_out_4;
                sbox_dout_aes_256_clk_26[23:16]   = AES_256_out_5;
                sbox_dout_aes_256_clk_26[15:8]    = AES_256_out_6;
                sbox_dout_aes_256_clk_26[7:0]     = AES_256_out_7;
                sbox_dout_aes_256_clk_26[127:120] = AES_256_out_12;
                sbox_dout_aes_256_clk_26[119:112] = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_26 = sbox_dout_aes_256_clk_26;
        endcase
    end else begin
        sbox_dout_aes_256_clk_26 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_26 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_26 = 32'h0;
        case (clk_cnt_all)
            6'h26: begin
                sbox_kout_aes_256_clk_26[31:24]   = AES_256_out_8;
                sbox_kout_aes_256_clk_26[23:16]   = AES_256_out_9;
                sbox_kout_aes_256_clk_26[15:8]    = AES_256_out_10;
                sbox_kout_aes_256_clk_26[7:0]     = AES_256_out_11;
            end
            default: sbox_kout_aes_256_clk_26 = sbox_kout_aes_256_clk_26;
        endcase
    end else begin
        sbox_kout_aes_256_clk_26 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_dout_aes_256_clk_27 = 128'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_dout_aes_256_clk_27 = 128'h0;
        case (clk_cnt_all)
            6'h27: begin
                sbox_dout_aes_256_clk_27[111:104] = AES_256_out_0;
                sbox_dout_aes_256_clk_27[103:96]  = AES_256_out_1;
                sbox_dout_aes_256_clk_27[95:88]   = AES_256_out_2;
                sbox_dout_aes_256_clk_27[87:80]   = AES_256_out_3;
                sbox_dout_aes_256_clk_27[79:72]   = AES_256_out_4;
                sbox_dout_aes_256_clk_27[71:64]   = AES_256_out_5;
                sbox_dout_aes_256_clk_27[63:56]   = AES_256_out_6;
                sbox_dout_aes_256_clk_27[55:48]   = AES_256_out_7;
                sbox_dout_aes_256_clk_27[47:40]   = AES_256_out_8;
                sbox_dout_aes_256_clk_27[39:32]   = AES_256_out_9;
                sbox_dout_aes_256_clk_27[31:24]   = AES_256_out_10;
                sbox_dout_aes_256_clk_27[23:16]   = AES_256_out_11;
                sbox_dout_aes_256_clk_27[15:8]    = AES_256_out_12;
                sbox_dout_aes_256_clk_27[7:0]     = AES_256_out_13;
            end
            default: sbox_dout_aes_256_clk_27 = sbox_dout_aes_256_clk_27;
        endcase
    end else begin
        sbox_dout_aes_256_clk_27 = 128'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_0 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_0 = 32'h0;
    end else begin
        BK_0_round_0 = 32'h0;
        case (clk_cnt_all)
            6'h0: begin
                BK_0_round_0[31:24] = SM4_out_0;
                BK_0_round_0[23:16] = SM4_out_1;
                BK_0_round_0[15:8]  = SM4_out_2;
                BK_0_round_0[7:0]   = SM4_out_3;
            end
            default: BK_0_round_0 = BK_0_round_0;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_0 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_0 = 32'h0;
    end else begin
        B_0_round_0 = 32'h0;
        case (clk_cnt_all)
            6'h0: begin
                B_0_round_0[31:24]  = SM4_out_4;
                B_0_round_0[23:16]  = SM4_out_5;
                B_0_round_0[15:8]   = SM4_out_6;
                B_0_round_0[7:0]    = SM4_out_7;
            end
            default: B_0_round_0 = B_0_round_0;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_1 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_1 = 32'h0;
    end else begin
        BK_1_round_1 = 32'h0;
        case (clk_cnt_all)
            6'h0: begin
                BK_1_round_1[31:24] = SM4_out_8;
                BK_1_round_1[23:16] = SM4_out_9;
                BK_1_round_1[15:8]  = SM4_out_10;
                BK_1_round_1[7:0]   = SM4_out_11;
            end
            default: BK_1_round_1 = BK_1_round_1;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_1 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_1 = 32'h0;
    end else begin
        B_1_round_1 = 32'h0;
        case (clk_cnt_all)
            6'h0: begin
                B_1_round_1[31:24]  = SM4_out_12;
            end
            6'h1: begin
                B_1_round_1[23:16]  = SM4_out_0;
                B_1_round_1[15:8]   = SM4_out_1;
                B_1_round_1[7:0]    = SM4_out_2;
            end
            default: B_1_round_1 = B_1_round_1;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_2 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_2 = 32'h0;
    end else begin
        BK_0_round_2 = 32'h0;
        case (clk_cnt_all)
            6'h1: begin
                BK_0_round_2[31:24] = SM4_out_3;
                BK_0_round_2[23:16] = SM4_out_4;
                BK_0_round_2[15:8]  = SM4_out_5;
                BK_0_round_2[7:0]   = SM4_out_6;
            end
            default: BK_0_round_2 = BK_0_round_2;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_2 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_2 = 32'h0;
    end else begin
        B_0_round_2 = 32'h0;
        case (clk_cnt_all)
            6'h1: begin
                B_0_round_2[31:24]  = SM4_out_7;
                B_0_round_2[23:16]  = SM4_out_8;
                B_0_round_2[15:8]   = SM4_out_9;
                B_0_round_2[7:0]    = SM4_out_10;
            end
            default: B_0_round_2 = B_0_round_2;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_3 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_3 = 32'h0;
    end else begin
        BK_1_round_3 = 32'h0;
        case (clk_cnt_all)
            6'h1: begin
                BK_1_round_3[31:24] = SM4_out_11;
                BK_1_round_3[23:16] = SM4_out_12;
            end
            6'h2: begin
                BK_1_round_3[15:8]  = SM4_out_0;
                BK_1_round_3[7:0]   = SM4_out_1;
            end
            default: BK_1_round_3 = BK_1_round_3;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_3 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_3 = 32'h0;
    end else begin
        B_1_round_3 = 32'h0;
        case (clk_cnt_all)
            6'h2: begin
                B_1_round_3[31:24]  = SM4_out_2;
                B_1_round_3[23:16]  = SM4_out_3;
                B_1_round_3[15:8]   = SM4_out_4;
                B_1_round_3[7:0]    = SM4_out_5;
            end
            default: B_1_round_3 = B_1_round_3;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_4 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_4 = 32'h0;
    end else begin
        BK_0_round_4 = 32'h0;
        case (clk_cnt_all)
            6'h2: begin
                BK_0_round_4[31:24] = SM4_out_6;
                BK_0_round_4[23:16] = SM4_out_7;
                BK_0_round_4[15:8]  = SM4_out_8;
                BK_0_round_4[7:0]   = SM4_out_9;
            end
            default: BK_0_round_4 = BK_0_round_4;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_4 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_4 = 32'h0;
    end else begin
        B_0_round_4 = 32'h0;
        case (clk_cnt_all)
            6'h2: begin
                B_0_round_4[31:24]  = SM4_out_10;
                B_0_round_4[23:16]  = SM4_out_11;
                B_0_round_4[15:8]   = SM4_out_12;
            end
            6'h3: begin
                B_0_round_4[7:0]    = SM4_out_0;
            end
            default: B_0_round_4 = B_0_round_4;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_5 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_5 = 32'h0;
    end else begin
        BK_1_round_5 = 32'h0;
        case (clk_cnt_all)
            6'h3: begin
                BK_1_round_5[31:24] = SM4_out_1;
                BK_1_round_5[23:16] = SM4_out_2;
                BK_1_round_5[15:8]  = SM4_out_3;
                BK_1_round_5[7:0]   = SM4_out_4;
            end
            default: BK_1_round_5 = BK_1_round_5;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_5 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_5 = 32'h0;
    end else begin
        B_1_round_5 = 32'h0;
        case (clk_cnt_all)
            6'h3: begin
                B_1_round_5[31:24]  = SM4_out_5;
                B_1_round_5[23:16]  = SM4_out_6;
                B_1_round_5[15:8]   = SM4_out_7;
                B_1_round_5[7:0]    = SM4_out_8;
            end
            default: B_1_round_5 = B_1_round_5;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_6 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_6 = 32'h0;
    end else begin
        BK_0_round_6 = 32'h0;
        case (clk_cnt_all)
            6'h3: begin
                BK_0_round_6[31:24] = SM4_out_9;
                BK_0_round_6[23:16] = SM4_out_10;
                BK_0_round_6[15:8]  = SM4_out_11;
                BK_0_round_6[7:0]   = SM4_out_12;
            end
            default: BK_0_round_6 = BK_0_round_6;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_6 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_6 = 32'h0;
    end else begin
        B_0_round_6 = 32'h0;
        case (clk_cnt_all)
            6'h4: begin
                B_0_round_6[31:24]  = SM4_out_0;
                B_0_round_6[23:16]  = SM4_out_1;
                B_0_round_6[15:8]   = SM4_out_2;
                B_0_round_6[7:0]    = SM4_out_3;
            end
            default: B_0_round_6 = B_0_round_6;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_7 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_7 = 32'h0;
    end else begin
        BK_1_round_7 = 32'h0;
        case (clk_cnt_all)
            6'h4: begin
                BK_1_round_7[31:24] = SM4_out_4;
                BK_1_round_7[23:16] = SM4_out_5;
                BK_1_round_7[15:8]  = SM4_out_6;
                BK_1_round_7[7:0]   = SM4_out_7;
            end
            default: BK_1_round_7 = BK_1_round_7;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_7 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_7 = 32'h0;
    end else begin
        B_1_round_7 = 32'h0;
        case (clk_cnt_all)
            6'h4: begin
                B_1_round_7[31:24]  = SM4_out_8;
                B_1_round_7[23:16]  = SM4_out_9;
                B_1_round_7[15:8]   = SM4_out_10;
                B_1_round_7[7:0]    = SM4_out_11;
            end
            default: B_1_round_7 = B_1_round_7;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_8 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_8 = 32'h0;
    end else begin
        BK_0_round_8 = 32'h0;
        case (clk_cnt_all)
            6'h4: begin
                BK_0_round_8[31:24] = SM4_out_12;
            end
            6'h5: begin
                BK_0_round_8[23:16] = SM4_out_0;
                BK_0_round_8[15:8]  = SM4_out_1;
                BK_0_round_8[7:0]   = SM4_out_2;
            end
            default: BK_0_round_8 = BK_0_round_8;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_8 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_8 = 32'h0;
    end else begin
        B_0_round_8 = 32'h0;
        case (clk_cnt_all)
            6'h5: begin
                B_0_round_8[31:24]  = SM4_out_3;
                B_0_round_8[23:16]  = SM4_out_4;
                B_0_round_8[15:8]   = SM4_out_5;
                B_0_round_8[7:0]    = SM4_out_6;
            end
            default: B_0_round_8 = B_0_round_8;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_9 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_9 = 32'h0;
    end else begin
        BK_1_round_9 = 32'h0;
        case (clk_cnt_all)
            6'h5: begin
                BK_1_round_9[31:24] = SM4_out_7;
                BK_1_round_9[23:16] = SM4_out_8;
                BK_1_round_9[15:8]  = SM4_out_9;
                BK_1_round_9[7:0]   = SM4_out_10;
            end
            default: BK_1_round_9 = BK_1_round_9;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_9 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_9 = 32'h0;
    end else begin
        B_1_round_9 = 32'h0;
        case (clk_cnt_all)
            6'h5: begin
                B_1_round_9[31:24]  = SM4_out_11;
                B_1_round_9[23:16]  = SM4_out_12;
            end
            6'h6: begin
                B_1_round_9[15:8]   = SM4_out_0;
                B_1_round_9[7:0]    = SM4_out_1;
            end
            default: B_1_round_9 = B_1_round_9;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_10 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_10 = 32'h0;
    end else begin
        BK_0_round_10 = 32'h0;
        case (clk_cnt_all)
            6'h6: begin
                BK_0_round_10[31:24]= SM4_out_2;
                BK_0_round_10[23:16]= SM4_out_3;
                BK_0_round_10[15:8] = SM4_out_4;
                BK_0_round_10[7:0]  = SM4_out_5;
            end
            default: BK_0_round_10 = BK_0_round_10;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_10 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_10 = 32'h0;
    end else begin
        B_0_round_10 = 32'h0;
        case (clk_cnt_all)
            6'h6: begin
                B_0_round_10[31:24] = SM4_out_6;
                B_0_round_10[23:16] = SM4_out_7;
                B_0_round_10[15:8]  = SM4_out_8;
                B_0_round_10[7:0]   = SM4_out_9;
            end
            default: B_0_round_10 = B_0_round_10;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_11 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_11 = 32'h0;
    end else begin
        BK_1_round_11 = 32'h0;
        case (clk_cnt_all)
            6'h6: begin
                BK_1_round_11[31:24]= SM4_out_10;
                BK_1_round_11[23:16]= SM4_out_11;
                BK_1_round_11[15:8] = SM4_out_12;
            end
            6'h7: begin
                BK_1_round_11[7:0]  = SM4_out_0;
            end
            default: BK_1_round_11 = BK_1_round_11;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_11 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_11 = 32'h0;
    end else begin
        B_1_round_11 = 32'h0;
        case (clk_cnt_all)
            6'h7: begin
                B_1_round_11[31:24] = SM4_out_1;
                B_1_round_11[23:16] = SM4_out_2;
                B_1_round_11[15:8]  = SM4_out_3;
                B_1_round_11[7:0]   = SM4_out_4;
            end
            default: B_1_round_11 = B_1_round_11;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_12 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_12 = 32'h0;
    end else begin
        BK_0_round_12 = 32'h0;
        case (clk_cnt_all)
            6'h7: begin
                BK_0_round_12[31:24]= SM4_out_5;
                BK_0_round_12[23:16]= SM4_out_6;
                BK_0_round_12[15:8] = SM4_out_7;
                BK_0_round_12[7:0]  = SM4_out_8;
            end
            default: BK_0_round_12 = BK_0_round_12;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_12 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_12 = 32'h0;
    end else begin
        B_0_round_12 = 32'h0;
        case (clk_cnt_all)
            6'h7: begin
                B_0_round_12[31:24] = SM4_out_9;
                B_0_round_12[23:16] = SM4_out_10;
                B_0_round_12[15:8]  = SM4_out_11;
                B_0_round_12[7:0]   = SM4_out_12;
            end
            default: B_0_round_12 = B_0_round_12;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_13 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_13 = 32'h0;
    end else begin
        BK_1_round_13 = 32'h0;
        case (clk_cnt_all)
            6'h8: begin
                BK_1_round_13[31:24]= SM4_out_0;
                BK_1_round_13[23:16]= SM4_out_1;
                BK_1_round_13[15:8] = SM4_out_2;
                BK_1_round_13[7:0]  = SM4_out_3;
            end
            default: BK_1_round_13 = BK_1_round_13;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_13 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_13 = 32'h0;
    end else begin
        B_1_round_13 = 32'h0;
        case (clk_cnt_all)
            6'h8: begin
                B_1_round_13[31:24] = SM4_out_4;
                B_1_round_13[23:16] = SM4_out_5;
                B_1_round_13[15:8]  = SM4_out_6;
                B_1_round_13[7:0]   = SM4_out_7;
            end
            default: B_1_round_13 = B_1_round_13;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_14 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_14 = 32'h0;
    end else begin
        BK_0_round_14 = 32'h0;
        case (clk_cnt_all)
            6'h8: begin
                BK_0_round_14[31:24]= SM4_out_8;
                BK_0_round_14[23:16]= SM4_out_9;
                BK_0_round_14[15:8] = SM4_out_10;
                BK_0_round_14[7:0]  = SM4_out_11;
            end
            default: BK_0_round_14 = BK_0_round_14;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_14 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_14 = 32'h0;
    end else begin
        B_0_round_14 = 32'h0;
        case (clk_cnt_all)
            6'h8: begin
                B_0_round_14[31:24] = SM4_out_12;
            end
            6'h9: begin
                B_0_round_14[23:16] = SM4_out_0;
                B_0_round_14[15:8]  = SM4_out_1;
                B_0_round_14[7:0]   = SM4_out_2;
            end
            default: B_0_round_14 = B_0_round_14;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_15 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_15 = 32'h0;
    end else begin
        BK_1_round_15 = 32'h0;
        case (clk_cnt_all)
            6'h9: begin
                BK_1_round_15[31:24]= SM4_out_3;
                BK_1_round_15[23:16]= SM4_out_4;
                BK_1_round_15[15:8] = SM4_out_5;
                BK_1_round_15[7:0]  = SM4_out_6;
            end
            default: BK_1_round_15 = BK_1_round_15;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_15 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_15 = 32'h0;
    end else begin
        B_1_round_15 = 32'h0;
        case (clk_cnt_all)
            6'h9: begin
                B_1_round_15[31:24] = SM4_out_7;
                B_1_round_15[23:16] = SM4_out_8;
                B_1_round_15[15:8]  = SM4_out_9;
                B_1_round_15[7:0]   = SM4_out_10;
            end
            default: B_1_round_15 = B_1_round_15;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_16 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_16 = 32'h0;
    end else begin
        BK_0_round_16 = 32'h0;
        case (clk_cnt_all)
            6'h9: begin
                BK_0_round_16[31:24]= SM4_out_11;
                BK_0_round_16[23:16]= SM4_out_12;
            end
            6'ha: begin
                BK_0_round_16[15:8] = SM4_out_0;
                BK_0_round_16[7:0]  = SM4_out_1;
            end
            default: BK_0_round_16 = BK_0_round_16;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_16 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_16 = 32'h0;
    end else begin
        B_0_round_16 = 32'h0;
        case (clk_cnt_all)
            6'ha: begin
                B_0_round_16[31:24] = SM4_out_2;
                B_0_round_16[23:16] = SM4_out_3;
                B_0_round_16[15:8]  = SM4_out_4;
                B_0_round_16[7:0]   = SM4_out_5;
            end
            default: B_0_round_16 = B_0_round_16;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_17 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_17 = 32'h0;
    end else begin
        BK_1_round_17 = 32'h0;
        case (clk_cnt_all)
            6'ha: begin
                BK_1_round_17[31:24]= SM4_out_6;
                BK_1_round_17[23:16]= SM4_out_7;
                BK_1_round_17[15:8] = SM4_out_8;
                BK_1_round_17[7:0]  = SM4_out_9;
            end
            default: BK_1_round_17 = BK_1_round_17;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_17 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_17 = 32'h0;
    end else begin
        B_1_round_17 = 32'h0;
        case (clk_cnt_all)
            6'ha: begin
                B_1_round_17[31:24] = SM4_out_10;
                B_1_round_17[23:16] = SM4_out_11;
                B_1_round_17[15:8]  = SM4_out_12;
            end
            6'hb: begin
                B_1_round_17[7:0]   = SM4_out_0;
            end
            default: B_1_round_17 = B_1_round_17;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_18 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_18 = 32'h0;
    end else begin
        BK_0_round_18 = 32'h0;
        case (clk_cnt_all)
            6'hb: begin
                BK_0_round_18[31:24]= SM4_out_1;
                BK_0_round_18[23:16]= SM4_out_2;
                BK_0_round_18[15:8] = SM4_out_3;
                BK_0_round_18[7:0]  = SM4_out_4;
            end
            default: BK_0_round_18 = BK_0_round_18;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_18 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_18 = 32'h0;
    end else begin
        B_0_round_18 = 32'h0;
        case (clk_cnt_all)
            6'hb: begin
                B_0_round_18[31:24] = SM4_out_5;
                B_0_round_18[23:16] = SM4_out_6;
                B_0_round_18[15:8]  = SM4_out_7;
                B_0_round_18[7:0]   = SM4_out_8;
            end
            default: B_0_round_18 = B_0_round_18;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_19 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_19 = 32'h0;
    end else begin
        BK_1_round_19 = 32'h0;
        case (clk_cnt_all)
            6'hb: begin
                BK_1_round_19[31:24]= SM4_out_9;
                BK_1_round_19[23:16]= SM4_out_10;
                BK_1_round_19[15:8] = SM4_out_11;
                BK_1_round_19[7:0]  = SM4_out_12;
            end
            default: BK_1_round_19 = BK_1_round_19;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_19 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_19 = 32'h0;
    end else begin
        B_1_round_19 = 32'h0;
        case (clk_cnt_all)
            6'hc: begin
                B_1_round_19[31:24] = SM4_out_0;
                B_1_round_19[23:16] = SM4_out_1;
                B_1_round_19[15:8]  = SM4_out_2;
                B_1_round_19[7:0]   = SM4_out_3;
            end
            default: B_1_round_19 = B_1_round_19;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_20 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_20 = 32'h0;
    end else begin
        BK_0_round_20 = 32'h0;
        case (clk_cnt_all)
            6'hc: begin
                BK_0_round_20[31:24]= SM4_out_4;
                BK_0_round_20[23:16]= SM4_out_5;
                BK_0_round_20[15:8] = SM4_out_6;
                BK_0_round_20[7:0]  = SM4_out_7;
            end
            default: BK_0_round_20 = BK_0_round_20;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_20 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_20 = 32'h0;
    end else begin
        B_0_round_20 = 32'h0;
        case (clk_cnt_all)
            6'hc: begin
                B_0_round_20[31:24] = SM4_out_8;
                B_0_round_20[23:16] = SM4_out_9;
                B_0_round_20[15:8]  = SM4_out_10;
                B_0_round_20[7:0]   = SM4_out_11;
            end
            default: B_0_round_20 = B_0_round_20;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_21 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_21 = 32'h0;
    end else begin
        BK_1_round_21 = 32'h0;
        case (clk_cnt_all)
            6'hc: begin
                BK_1_round_21[31:24]= SM4_out_12;
            end
            6'hd: begin
                BK_1_round_21[23:16]= SM4_out_0;
                BK_1_round_21[15:8] = SM4_out_1;
                BK_1_round_21[7:0]  = SM4_out_2;
            end
            default: BK_1_round_21 = BK_1_round_21;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_21 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_21 = 32'h0;
    end else begin
        B_1_round_21 = 32'h0;
        case (clk_cnt_all)
            6'hd: begin
                B_1_round_21[31:24] = SM4_out_3;
                B_1_round_21[23:16] = SM4_out_4;
                B_1_round_21[15:8]  = SM4_out_5;
                B_1_round_21[7:0]   = SM4_out_6;
            end
            default: B_1_round_21 = B_1_round_21;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_22 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_22 = 32'h0;
    end else begin
        BK_0_round_22 = 32'h0;
        case (clk_cnt_all)
            6'hd: begin
                BK_0_round_22[31:24]= SM4_out_7;
                BK_0_round_22[23:16]= SM4_out_8;
                BK_0_round_22[15:8] = SM4_out_9;
                BK_0_round_22[7:0]  = SM4_out_10;
            end
            default: BK_0_round_22 = BK_0_round_22;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_22 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_22 = 32'h0;
    end else begin
        B_0_round_22 = 32'h0;
        case (clk_cnt_all)
            6'hd: begin
                B_0_round_22[31:24] = SM4_out_11;
                B_0_round_22[23:16] = SM4_out_12;
            end
            6'he: begin
                B_0_round_22[15:8]  = SM4_out_0;
                B_0_round_22[7:0]   = SM4_out_1;
            end
            default: B_0_round_22 = B_0_round_22;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_23 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_23 = 32'h0;
    end else begin
        BK_1_round_23 = 32'h0;
        case (clk_cnt_all)
            6'he: begin
                BK_1_round_23[31:24]= SM4_out_2;
                BK_1_round_23[23:16]= SM4_out_3;
                BK_1_round_23[15:8] = SM4_out_4;
                BK_1_round_23[7:0]  = SM4_out_5;
            end
            default: BK_1_round_23 = BK_1_round_23;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_23 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_23 = 32'h0;
    end else begin
        B_1_round_23 = 32'h0;
        case (clk_cnt_all)
            6'he: begin
                B_1_round_23[31:24] = SM4_out_6;
                B_1_round_23[23:16] = SM4_out_7;
                B_1_round_23[15:8]  = SM4_out_8;
                B_1_round_23[7:0]   = SM4_out_9;
            end
            default: B_1_round_23 = B_1_round_23;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_24 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_24 = 32'h0;
    end else begin
        BK_0_round_24 = 32'h0;
        case (clk_cnt_all)
            6'he: begin
                BK_0_round_24[31:24]= SM4_out_10;
                BK_0_round_24[23:16]= SM4_out_11;
                BK_0_round_24[15:8] = SM4_out_12;
            end
            6'hf: begin
                BK_0_round_24[7:0]  = SM4_out_0;
            end
            default: BK_0_round_24 = BK_0_round_24;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_24 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_24 = 32'h0;
    end else begin
        B_0_round_24 = 32'h0;
        case (clk_cnt_all)
            6'hf: begin
                B_0_round_24[31:24] = SM4_out_1;
                B_0_round_24[23:16] = SM4_out_2;
                B_0_round_24[15:8]  = SM4_out_3;
                B_0_round_24[7:0]   = SM4_out_4;
            end
            default: B_0_round_24 = B_0_round_24;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_25 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_25 = 32'h0;
    end else begin
        BK_1_round_25 = 32'h0;
        case (clk_cnt_all)
            6'hf: begin
                BK_1_round_25[31:24]= SM4_out_5;
                BK_1_round_25[23:16]= SM4_out_6;
                BK_1_round_25[15:8] = SM4_out_7;
                BK_1_round_25[7:0]  = SM4_out_8;
            end
            default: BK_1_round_25 = BK_1_round_25;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_25 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_25 = 32'h0;
    end else begin
        B_1_round_25 = 32'h0;
        case (clk_cnt_all)
            6'hf: begin
                B_1_round_25[31:24] = SM4_out_9;
                B_1_round_25[23:16] = SM4_out_10;
                B_1_round_25[15:8]  = SM4_out_11;
                B_1_round_25[7:0]   = SM4_out_12;
            end
            default: B_1_round_25 = B_1_round_25;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_26 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_26 = 32'h0;
    end else begin
        BK_0_round_26 = 32'h0;
        case (clk_cnt_all)
            6'h10: begin
                BK_0_round_26[31:24]= SM4_out_0;
                BK_0_round_26[23:16]= SM4_out_1;
                BK_0_round_26[15:8] = SM4_out_2;
                BK_0_round_26[7:0]  = SM4_out_3;
            end
            default: BK_0_round_26 = BK_0_round_26;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_26 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_26 = 32'h0;
    end else begin
        B_0_round_26 = 32'h0;
        case (clk_cnt_all)
            6'h10: begin
                B_0_round_26[31:24] = SM4_out_4;
                B_0_round_26[23:16] = SM4_out_5;
                B_0_round_26[15:8]  = SM4_out_6;
                B_0_round_26[7:0]   = SM4_out_7;
            end
            default: B_0_round_26 = B_0_round_26;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_27 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_27 = 32'h0;
    end else begin
        BK_1_round_27 = 32'h0;
        case (clk_cnt_all)
            6'h10: begin
                BK_1_round_27[31:24]= SM4_out_8;
                BK_1_round_27[23:16]= SM4_out_9;
                BK_1_round_27[15:8] = SM4_out_10;
                BK_1_round_27[7:0]  = SM4_out_11;
            end
            default: BK_1_round_27 = BK_1_round_27;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_27 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_27 = 32'h0;
    end else begin
        B_1_round_27 = 32'h0;
        case (clk_cnt_all)
            6'h10: begin
                B_1_round_27[31:24] = SM4_out_12;
            end
            6'h11: begin
                B_1_round_27[23:16] = SM4_out_0;
                B_1_round_27[15:8]  = SM4_out_1;
                B_1_round_27[7:0]   = SM4_out_2;
            end
            default: B_1_round_27 = B_1_round_27;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_28 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_28 = 32'h0;
    end else begin
        BK_0_round_28 = 32'h0;
        case (clk_cnt_all)
            6'h11: begin
                BK_0_round_28[31:24]= SM4_out_3;
                BK_0_round_28[23:16]= SM4_out_4;
                BK_0_round_28[15:8] = SM4_out_5;
                BK_0_round_28[7:0]  = SM4_out_6;
            end
            default: BK_0_round_28 = BK_0_round_28;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_28 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_28 = 32'h0;
    end else begin
        B_0_round_28 = 32'h0;
        case (clk_cnt_all)
            6'h11: begin
                B_0_round_28[31:24] = SM4_out_7;
                B_0_round_28[23:16] = SM4_out_8;
                B_0_round_28[15:8]  = SM4_out_9;
                B_0_round_28[7:0]   = SM4_out_10;
            end
            default: B_0_round_28 = B_0_round_28;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_29 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_29 = 32'h0;
    end else begin
        BK_1_round_29 = 32'h0;
        case (clk_cnt_all)
            6'h11: begin
                BK_1_round_29[31:24]= SM4_out_11;
                BK_1_round_29[23:16]= SM4_out_12;
            end
            6'h12: begin
                BK_1_round_29[15:8] = SM4_out_0;
                BK_1_round_29[7:0]  = SM4_out_1;
            end
            default: BK_1_round_29 = BK_1_round_29;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_29 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_29 = 32'h0;
    end else begin
        B_1_round_29 = 32'h0;
        case (clk_cnt_all)
            6'h12: begin
                B_1_round_29[31:24] = SM4_out_2;
                B_1_round_29[23:16] = SM4_out_3;
                B_1_round_29[15:8]  = SM4_out_4;
                B_1_round_29[7:0]   = SM4_out_5;
            end
            default: B_1_round_29 = B_1_round_29;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_30 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_30 = 32'h0;
    end else begin
        BK_0_round_30 = 32'h0;
        case (clk_cnt_all)
            6'h12: begin
                BK_0_round_30[31:24]= SM4_out_6;
                BK_0_round_30[23:16]= SM4_out_7;
                BK_0_round_30[15:8] = SM4_out_8;
                BK_0_round_30[7:0]  = SM4_out_9;
            end
            default: BK_0_round_30 = BK_0_round_30;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_30 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_30 = 32'h0;
    end else begin
        B_0_round_30 = 32'h0;
        case (clk_cnt_all)
            6'h12: begin
                B_0_round_30[31:24] = SM4_out_10;
                B_0_round_30[23:16] = SM4_out_11;
                B_0_round_30[15:8]  = SM4_out_12;
            end
            6'h13: begin
                B_0_round_30[7:0]   = SM4_out_0;
            end
            default: B_0_round_30 = B_0_round_30;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_31 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_31 = 32'h0;
    end else begin
        BK_1_round_31 = 32'h0;
        case (clk_cnt_all)
            6'h13: begin
                BK_1_round_31[31:24]= SM4_out_1;
                BK_1_round_31[23:16]= SM4_out_2;
                BK_1_round_31[15:8] = SM4_out_3;
                BK_1_round_31[7:0]  = SM4_out_4;
            end
            default: BK_1_round_31 = BK_1_round_31;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_31 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_31 = 32'h0;
    end else begin
        B_1_round_31 = 32'h0;
        case (clk_cnt_all)
            6'h13: begin
                B_1_round_31[31:24] = SM4_out_5;
                B_1_round_31[23:16] = SM4_out_6;
                B_1_round_31[15:8]  = SM4_out_7;
                B_1_round_31[7:0]   = SM4_out_8;
            end
            default: B_1_round_31 = B_1_round_31;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_32 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_32 = 32'h0;
    end else begin
        BK_0_round_32 = 32'h0;
        case (clk_cnt_all)
            6'h14: begin
                BK_0_round_32[31:24]= SM4_out_0;
                BK_0_round_32[23:16]= SM4_out_1;
                BK_0_round_32[15:8] = SM4_out_2;
                BK_0_round_32[7:0]  = SM4_out_3;
            end
            default: BK_0_round_32 = BK_0_round_32;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_32 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_32 = 32'h0;
    end else begin
        B_0_round_32 = 32'h0;
        case (clk_cnt_all)
            6'h14: begin
                B_0_round_32[31:24] = SM4_out_4;
                B_0_round_32[23:16] = SM4_out_5;
                B_0_round_32[15:8]  = SM4_out_6;
                B_0_round_32[7:0]   = SM4_out_7;
            end
            default: B_0_round_32 = B_0_round_32;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_33 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_33 = 32'h0;
    end else begin
        BK_1_round_33 = 32'h0;
        case (clk_cnt_all)
            6'h14: begin
                BK_1_round_33[31:24]= SM4_out_8;
                BK_1_round_33[23:16]= SM4_out_9;
                BK_1_round_33[15:8] = SM4_out_10;
                BK_1_round_33[7:0]  = SM4_out_11;
            end
            default: BK_1_round_33 = BK_1_round_33;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_33 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_33 = 32'h0;
    end else begin
        B_1_round_33 = 32'h0;
        case (clk_cnt_all)
            6'h14: begin
                B_1_round_33[31:24] = SM4_out_12;
            end
            6'h15: begin
                B_1_round_33[23:16] = SM4_out_0;
                B_1_round_33[15:8]  = SM4_out_1;
                B_1_round_33[7:0]   = SM4_out_2;
            end
            default: B_1_round_33 = B_1_round_33;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_34 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_34 = 32'h0;
    end else begin
        BK_0_round_34 = 32'h0;
        case (clk_cnt_all)
            6'h15: begin
                BK_0_round_34[31:24]= SM4_out_3;
                BK_0_round_34[23:16]= SM4_out_4;
                BK_0_round_34[15:8] = SM4_out_5;
                BK_0_round_34[7:0]  = SM4_out_6;
            end
            default: BK_0_round_34 = BK_0_round_34;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_34 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_34 = 32'h0;
    end else begin
        B_0_round_34 = 32'h0;
        case (clk_cnt_all)
            6'h15: begin
                B_0_round_34[31:24] = SM4_out_7;
                B_0_round_34[23:16] = SM4_out_8;
                B_0_round_34[15:8]  = SM4_out_9;
                B_0_round_34[7:0]   = SM4_out_10;
            end
            default: B_0_round_34 = B_0_round_34;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_35 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_35 = 32'h0;
    end else begin
        BK_1_round_35 = 32'h0;
        case (clk_cnt_all)
            6'h15: begin
                BK_1_round_35[31:24]= SM4_out_11;
                BK_1_round_35[23:16]= SM4_out_12;
            end
            6'h16: begin
                BK_1_round_35[15:8] = SM4_out_0;
                BK_1_round_35[7:0]  = SM4_out_1;
            end
            default: BK_1_round_35 = BK_1_round_35;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_35 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_35 = 32'h0;
    end else begin
        B_1_round_35 = 32'h0;
        case (clk_cnt_all)
            6'h16: begin
                B_1_round_35[31:24] = SM4_out_2;
                B_1_round_35[23:16] = SM4_out_3;
                B_1_round_35[15:8]  = SM4_out_4;
                B_1_round_35[7:0]   = SM4_out_5;
            end
            default: B_1_round_35 = B_1_round_35;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_36 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_36 = 32'h0;
    end else begin
        BK_0_round_36 = 32'h0;
        case (clk_cnt_all)
            6'h16: begin
                BK_0_round_36[31:24]= SM4_out_6;
                BK_0_round_36[23:16]= SM4_out_7;
                BK_0_round_36[15:8] = SM4_out_8;
                BK_0_round_36[7:0]  = SM4_out_9;
            end
            default: BK_0_round_36 = BK_0_round_36;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_36 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_36 = 32'h0;
    end else begin
        B_0_round_36 = 32'h0;
        case (clk_cnt_all)
            6'h16: begin
                B_0_round_36[31:24] = SM4_out_10;
                B_0_round_36[23:16] = SM4_out_11;
                B_0_round_36[15:8]  = SM4_out_12;
            end
            6'h17: begin
                B_0_round_36[7:0]   = SM4_out_0;
            end
            default: B_0_round_36 = B_0_round_36;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_37 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_37 = 32'h0;
    end else begin
        BK_1_round_37 = 32'h0;
        case (clk_cnt_all)
            6'h17: begin
                BK_1_round_37[31:24]= SM4_out_1;
                BK_1_round_37[23:16]= SM4_out_2;
                BK_1_round_37[15:8] = SM4_out_3;
                BK_1_round_37[7:0]  = SM4_out_4;
            end
            default: BK_1_round_37 = BK_1_round_37;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_37 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_37 = 32'h0;
    end else begin
        B_1_round_37 = 32'h0;
        case (clk_cnt_all)
            6'h17: begin
                B_1_round_37[31:24] = SM4_out_5;
                B_1_round_37[23:16] = SM4_out_6;
                B_1_round_37[15:8]  = SM4_out_7;
                B_1_round_37[7:0]   = SM4_out_8;
            end
            default: B_1_round_37 = B_1_round_37;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_38 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_38 = 32'h0;
    end else begin
        BK_0_round_38 = 32'h0;
        case (clk_cnt_all)
            6'h17: begin
                BK_0_round_38[31:24]= SM4_out_9;
                BK_0_round_38[23:16]= SM4_out_10;
                BK_0_round_38[15:8] = SM4_out_11;
                BK_0_round_38[7:0]  = SM4_out_12;
            end
            default: BK_0_round_38 = BK_0_round_38;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_38 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_38 = 32'h0;
    end else begin
        B_0_round_38 = 32'h0;
        case (clk_cnt_all)
            6'h18: begin
                B_0_round_38[31:24] = SM4_out_0;
                B_0_round_38[23:16] = SM4_out_1;
                B_0_round_38[15:8]  = SM4_out_2;
                B_0_round_38[7:0]   = SM4_out_3;
            end
            default: B_0_round_38 = B_0_round_38;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_39 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_39 = 32'h0;
    end else begin
        BK_1_round_39 = 32'h0;
        case (clk_cnt_all)
            6'h18: begin
                BK_1_round_39[31:24]= SM4_out_4;
                BK_1_round_39[23:16]= SM4_out_5;
                BK_1_round_39[15:8] = SM4_out_6;
                BK_1_round_39[7:0]  = SM4_out_7;
            end
            default: BK_1_round_39 = BK_1_round_39;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_39 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_39 = 32'h0;
    end else begin
        B_1_round_39 = 32'h0;
        case (clk_cnt_all)
            6'h18: begin
                B_1_round_39[31:24] = SM4_out_8;
                B_1_round_39[23:16] = SM4_out_9;
                B_1_round_39[15:8]  = SM4_out_10;
                B_1_round_39[7:0]   = SM4_out_11;
            end
            default: B_1_round_39 = B_1_round_39;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_40 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_40 = 32'h0;
    end else begin
        BK_0_round_40 = 32'h0;
        case (clk_cnt_all)
            6'h18: begin
                BK_0_round_40[31:24]= SM4_out_12;
            end
            6'h19: begin
                BK_0_round_40[23:16]= SM4_out_0;
                BK_0_round_40[15:8] = SM4_out_1;
                BK_0_round_40[7:0]  = SM4_out_2;
            end
            default: BK_0_round_40 = BK_0_round_40;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_40 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_40 = 32'h0;
    end else begin
        B_0_round_40 = 32'h0;
        case (clk_cnt_all)
            6'h19: begin
                B_0_round_40[31:24] = SM4_out_3;
                B_0_round_40[23:16] = SM4_out_4;
                B_0_round_40[15:8]  = SM4_out_5;
                B_0_round_40[7:0]   = SM4_out_6;
            end
            default: B_0_round_40 = B_0_round_40;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_41 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_41 = 32'h0;
    end else begin
        BK_1_round_41 = 32'h0;
        case (clk_cnt_all)
            6'h19: begin
                BK_1_round_41[31:24]= SM4_out_7;
                BK_1_round_41[23:16]= SM4_out_8;
                BK_1_round_41[15:8] = SM4_out_9;
                BK_1_round_41[7:0]  = SM4_out_10;
            end
            default: BK_1_round_41 = BK_1_round_41;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_41 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_41 = 32'h0;
    end else begin
        B_1_round_41 = 32'h0;
        case (clk_cnt_all)
            6'h19: begin
                B_1_round_41[31:24] = SM4_out_11;
                B_1_round_41[23:16] = SM4_out_12;
            end
            6'h1a: begin
                B_1_round_41[15:8]  = SM4_out_0;
                B_1_round_41[7:0]   = SM4_out_1;
            end
            default: B_1_round_41 = B_1_round_41;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_42 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_42 = 32'h0;
    end else begin
        BK_0_round_42 = 32'h0;
        case (clk_cnt_all)
            6'h1a: begin
                BK_0_round_42[31:24]= SM4_out_2;
                BK_0_round_42[23:16]= SM4_out_3;
                BK_0_round_42[15:8] = SM4_out_4;
                BK_0_round_42[7:0]  = SM4_out_5;
            end
            default: BK_0_round_42 = BK_0_round_42;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_42 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_42 = 32'h0;
    end else begin
        B_0_round_42 = 32'h0;
        case (clk_cnt_all)
            6'h1a: begin
                B_0_round_42[31:24] = SM4_out_6;
                B_0_round_42[23:16] = SM4_out_7;
                B_0_round_42[15:8]  = SM4_out_8;
                B_0_round_42[7:0]   = SM4_out_9;
            end
            default: B_0_round_42 = B_0_round_42;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_43 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_43 = 32'h0;
    end else begin
        BK_1_round_43 = 32'h0;
        case (clk_cnt_all)
            6'h1a: begin
                BK_1_round_43[31:24]= SM4_out_10;
                BK_1_round_43[23:16]= SM4_out_11;
                BK_1_round_43[15:8] = SM4_out_12;
            end
            6'h1b: begin
                BK_1_round_43[7:0]  = SM4_out_0;
            end
            default: BK_1_round_43 = BK_1_round_43;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_43 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_43 = 32'h0;
    end else begin
        B_1_round_43 = 32'h0;
        case (clk_cnt_all)
            6'h1b: begin
                B_1_round_43[31:24] = SM4_out_1;
                B_1_round_43[23:16] = SM4_out_2;
                B_1_round_43[15:8]  = SM4_out_3;
                B_1_round_43[7:0]   = SM4_out_4;
            end
            default: B_1_round_43 = B_1_round_43;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_44 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_44 = 32'h0;
    end else begin
        BK_0_round_44 = 32'h0;
        case (clk_cnt_all)
            6'h1b: begin
                BK_0_round_44[31:24]= SM4_out_5;
                BK_0_round_44[23:16]= SM4_out_6;
                BK_0_round_44[15:8] = SM4_out_7;
                BK_0_round_44[7:0]  = SM4_out_8;
            end
            default: BK_0_round_44 = BK_0_round_44;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_44 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_44 = 32'h0;
    end else begin
        B_0_round_44 = 32'h0;
        case (clk_cnt_all)
            6'h1b: begin
                B_0_round_44[31:24] = SM4_out_9;
                B_0_round_44[23:16] = SM4_out_10;
                B_0_round_44[15:8]  = SM4_out_11;
                B_0_round_44[7:0]   = SM4_out_12;
            end
            default: B_0_round_44 = B_0_round_44;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_45 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_45 = 32'h0;
    end else begin
        BK_1_round_45 = 32'h0;
        case (clk_cnt_all)
            6'h1c: begin
                BK_1_round_45[31:24]= SM4_out_0;
                BK_1_round_45[23:16]= SM4_out_1;
                BK_1_round_45[15:8] = SM4_out_2;
                BK_1_round_45[7:0]  = SM4_out_3;
            end
            default: BK_1_round_45 = BK_1_round_45;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_45 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_45 = 32'h0;
    end else begin
        B_1_round_45 = 32'h0;
        case (clk_cnt_all)
            6'h1c: begin
                B_1_round_45[31:24] = SM4_out_4;
                B_1_round_45[23:16] = SM4_out_5;
                B_1_round_45[15:8]  = SM4_out_6;
                B_1_round_45[7:0]   = SM4_out_7;
            end
            default: B_1_round_45 = B_1_round_45;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_46 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_46 = 32'h0;
    end else begin
        BK_0_round_46 = 32'h0;
        case (clk_cnt_all)
            6'h1c: begin
                BK_0_round_46[31:24]= SM4_out_8;
                BK_0_round_46[23:16]= SM4_out_9;
                BK_0_round_46[15:8] = SM4_out_10;
                BK_0_round_46[7:0]  = SM4_out_11;
            end
            default: BK_0_round_46 = BK_0_round_46;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_46 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_46 = 32'h0;
    end else begin
        B_0_round_46 = 32'h0;
        case (clk_cnt_all)
            6'h1c: begin
                B_0_round_46[31:24] = SM4_out_12;
            end
            6'h1d: begin
                B_0_round_46[23:16] = SM4_out_0;
                B_0_round_46[15:8]  = SM4_out_1;
                B_0_round_46[7:0]   = SM4_out_2;
            end
            default: B_0_round_46 = B_0_round_46;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_47 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_47 = 32'h0;
    end else begin
        BK_1_round_47 = 32'h0;
        case (clk_cnt_all)
            6'h1d: begin
                BK_1_round_47[31:24]= SM4_out_3;
                BK_1_round_47[23:16]= SM4_out_4;
                BK_1_round_47[15:8] = SM4_out_5;
                BK_1_round_47[7:0]  = SM4_out_6;
            end
            default: BK_1_round_47 = BK_1_round_47;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_47 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_47 = 32'h0;
    end else begin
        B_1_round_47 = 32'h0;
        case (clk_cnt_all)
            6'h1d: begin
                B_1_round_47[31:24] = SM4_out_7;
                B_1_round_47[23:16] = SM4_out_8;
                B_1_round_47[15:8]  = SM4_out_9;
                B_1_round_47[7:0]   = SM4_out_10;
            end
            default: B_1_round_47 = B_1_round_47;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_48 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_48 = 32'h0;
    end else begin
        BK_0_round_48 = 32'h0;
        case (clk_cnt_all)
            6'h1d: begin
                BK_0_round_48[31:24]= SM4_out_11;
                BK_0_round_48[23:16]= SM4_out_12;
            end
            6'h1e: begin
                BK_0_round_48[15:8] = SM4_out_0;
                BK_0_round_48[7:0]  = SM4_out_1;
            end
            default: BK_0_round_48 = BK_0_round_48;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_48 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_48 = 32'h0;
    end else begin
        B_0_round_48 = 32'h0;
        case (clk_cnt_all)
            6'h1e: begin
                B_0_round_48[31:24] = SM4_out_2;
                B_0_round_48[23:16] = SM4_out_3;
                B_0_round_48[15:8]  = SM4_out_4;
                B_0_round_48[7:0]   = SM4_out_5;
            end
            default: B_0_round_48 = B_0_round_48;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_49 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_49 = 32'h0;
    end else begin
        BK_1_round_49 = 32'h0;
        case (clk_cnt_all)
            6'h1e: begin
                BK_1_round_49[31:24]= SM4_out_6;
                BK_1_round_49[23:16]= SM4_out_7;
                BK_1_round_49[15:8] = SM4_out_8;
                BK_1_round_49[7:0]  = SM4_out_9;
            end
            default: BK_1_round_49 = BK_1_round_49;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_49 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_49 = 32'h0;
    end else begin
        B_1_round_49 = 32'h0;
        case (clk_cnt_all)
            6'h1e: begin
                B_1_round_49[31:24] = SM4_out_10;
                B_1_round_49[23:16] = SM4_out_11;
                B_1_round_49[15:8]  = SM4_out_12;
            end
            6'h1f: begin
                B_1_round_49[7:0]   = SM4_out_0;
            end
            default: B_1_round_49 = B_1_round_49;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_50 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_50 = 32'h0;
    end else begin
        BK_0_round_50 = 32'h0;
        case (clk_cnt_all)
            6'h1f: begin
                BK_0_round_50[31:24]= SM4_out_1;
                BK_0_round_50[23:16]= SM4_out_2;
                BK_0_round_50[15:8] = SM4_out_3;
                BK_0_round_50[7:0]  = SM4_out_4;
            end
            default: BK_0_round_50 = BK_0_round_50;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_50 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_50 = 32'h0;
    end else begin
        B_0_round_50 = 32'h0;
        case (clk_cnt_all)
            6'h1f: begin
                B_0_round_50[31:24] = SM4_out_5;
                B_0_round_50[23:16] = SM4_out_6;
                B_0_round_50[15:8]  = SM4_out_7;
                B_0_round_50[7:0]   = SM4_out_8;
            end
            default: B_0_round_50 = B_0_round_50;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_51 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_51 = 32'h0;
    end else begin
        BK_1_round_51 = 32'h0;
        case (clk_cnt_all)
            6'h1f: begin
                BK_1_round_51[31:24]= SM4_out_9;
                BK_1_round_51[23:16]= SM4_out_10;
                BK_1_round_51[15:8] = SM4_out_11;
                BK_1_round_51[7:0]  = SM4_out_12;
            end
            default: BK_1_round_51 = BK_1_round_51;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_51 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_51 = 32'h0;
    end else begin
        B_1_round_51 = 32'h0;
        case (clk_cnt_all)
            6'h20: begin
                B_1_round_51[31:24] = SM4_out_0;
                B_1_round_51[23:16] = SM4_out_1;
                B_1_round_51[15:8]  = SM4_out_2;
                B_1_round_51[7:0]   = SM4_out_3;
            end
            default: B_1_round_51 = B_1_round_51;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_52 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_52 = 32'h0;
    end else begin
        BK_0_round_52 = 32'h0;
        case (clk_cnt_all)
            6'h20: begin
                BK_0_round_52[31:24]= SM4_out_4;
                BK_0_round_52[23:16]= SM4_out_5;
                BK_0_round_52[15:8] = SM4_out_6;
                BK_0_round_52[7:0]  = SM4_out_7;
            end
            default: BK_0_round_52 = BK_0_round_52;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_52 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_52 = 32'h0;
    end else begin
        B_0_round_52 = 32'h0;
        case (clk_cnt_all)
            6'h20: begin
                B_0_round_52[31:24] = SM4_out_8;
                B_0_round_52[23:16] = SM4_out_9;
                B_0_round_52[15:8]  = SM4_out_10;
                B_0_round_52[7:0]   = SM4_out_11;
            end
            default: B_0_round_52 = B_0_round_52;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_53 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_53 = 32'h0;
    end else begin
        BK_1_round_53 = 32'h0;
        case (clk_cnt_all)
            6'h20: begin
                BK_1_round_53[31:24]= SM4_out_12;
            end
            6'h21: begin
                BK_1_round_53[23:16]= SM4_out_0;
                BK_1_round_53[15:8] = SM4_out_1;
                BK_1_round_53[7:0]  = SM4_out_2;
            end
            default: BK_1_round_53 = BK_1_round_53;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_53 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_53 = 32'h0;
    end else begin
        B_1_round_53 = 32'h0;
        case (clk_cnt_all)
            6'h21: begin
                B_1_round_53[31:24] = SM4_out_3;
                B_1_round_53[23:16] = SM4_out_4;
                B_1_round_53[15:8]  = SM4_out_5;
                B_1_round_53[7:0]   = SM4_out_6;
            end
            default: B_1_round_53 = B_1_round_53;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_54 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_54 = 32'h0;
    end else begin
        BK_0_round_54 = 32'h0;
        case (clk_cnt_all)
            6'h21: begin
                BK_0_round_54[31:24]= SM4_out_7;
                BK_0_round_54[23:16]= SM4_out_8;
                BK_0_round_54[15:8] = SM4_out_9;
                BK_0_round_54[7:0]  = SM4_out_10;
            end
            default: BK_0_round_54 = BK_0_round_54;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_54 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_54 = 32'h0;
    end else begin
        B_0_round_54 = 32'h0;
        case (clk_cnt_all)
            6'h21: begin
                B_0_round_54[31:24] = SM4_out_11;
                B_0_round_54[23:16] = SM4_out_12;
            end
            6'h22: begin
                B_0_round_54[15:8]  = SM4_out_0;
                B_0_round_54[7:0]   = SM4_out_1;
            end
            default: B_0_round_54 = B_0_round_54;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_55 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_55 = 32'h0;
    end else begin
        BK_1_round_55 = 32'h0;
        case (clk_cnt_all)
            6'h22: begin
                BK_1_round_55[31:24]= SM4_out_2;
                BK_1_round_55[23:16]= SM4_out_3;
                BK_1_round_55[15:8] = SM4_out_4;
                BK_1_round_55[7:0]  = SM4_out_5;
            end
            default: BK_1_round_55 = BK_1_round_55;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_55 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_55 = 32'h0;
    end else begin
        B_1_round_55 = 32'h0;
        case (clk_cnt_all)
            6'h22: begin
                B_1_round_55[31:24] = SM4_out_6;
                B_1_round_55[23:16] = SM4_out_7;
                B_1_round_55[15:8]  = SM4_out_8;
                B_1_round_55[7:0]   = SM4_out_9;
            end
            default: B_1_round_55 = B_1_round_55;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_56 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_56 = 32'h0;
    end else begin
        BK_0_round_56 = 32'h0;
        case (clk_cnt_all)
            6'h22: begin
                BK_0_round_56[31:24]= SM4_out_10;
                BK_0_round_56[23:16]= SM4_out_11;
                BK_0_round_56[15:8] = SM4_out_12;
            end
            6'h23: begin
                BK_0_round_56[7:0]  = SM4_out_0;
            end
            default: BK_0_round_56 = BK_0_round_56;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_56 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_56 = 32'h0;
    end else begin
        B_0_round_56 = 32'h0;
        case (clk_cnt_all)
            6'h23: begin
                B_0_round_56[31:24] = SM4_out_1;
                B_0_round_56[23:16] = SM4_out_2;
                B_0_round_56[15:8]  = SM4_out_3;
                B_0_round_56[7:0]   = SM4_out_4;
            end
            default: B_0_round_56 = B_0_round_56;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_57 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_57 = 32'h0;
    end else begin
        BK_1_round_57 = 32'h0;
        case (clk_cnt_all)
            6'h23: begin
                BK_1_round_57[31:24]= SM4_out_5;
                BK_1_round_57[23:16]= SM4_out_6;
                BK_1_round_57[15:8] = SM4_out_7;
                BK_1_round_57[7:0]  = SM4_out_8;
            end
            default: BK_1_round_57 = BK_1_round_57;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_57 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_57 = 32'h0;
    end else begin
        B_1_round_57 = 32'h0;
        case (clk_cnt_all)
            6'h23: begin
                B_1_round_57[31:24] = SM4_out_9;
                B_1_round_57[23:16] = SM4_out_10;
                B_1_round_57[15:8]  = SM4_out_11;
                B_1_round_57[7:0]   = SM4_out_12;
            end
            default: B_1_round_57 = B_1_round_57;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_58 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_58 = 32'h0;
    end else begin
        BK_0_round_58 = 32'h0;
        case (clk_cnt_all)
            6'h24: begin
                BK_0_round_58[31:24]= SM4_out_0;
                BK_0_round_58[23:16]= SM4_out_1;
                BK_0_round_58[15:8] = SM4_out_2;
                BK_0_round_58[7:0]  = SM4_out_3;
            end
            default: BK_0_round_58 = BK_0_round_58;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_58 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_58 = 32'h0;
    end else begin
        B_0_round_58 = 32'h0;
        case (clk_cnt_all)
            6'h24: begin
                B_0_round_58[31:24] = SM4_out_4;
                B_0_round_58[23:16] = SM4_out_5;
                B_0_round_58[15:8]  = SM4_out_6;
                B_0_round_58[7:0]   = SM4_out_7;
            end
            default: B_0_round_58 = B_0_round_58;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_59 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_59 = 32'h0;
    end else begin
        BK_1_round_59 = 32'h0;
        case (clk_cnt_all)
            6'h24: begin
                BK_1_round_59[31:24]= SM4_out_8;
                BK_1_round_59[23:16]= SM4_out_9;
                BK_1_round_59[15:8] = SM4_out_10;
                BK_1_round_59[7:0]  = SM4_out_11;
            end
            default: BK_1_round_59 = BK_1_round_59;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_59 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_59 = 32'h0;
    end else begin
        B_1_round_59 = 32'h0;
        case (clk_cnt_all)
            6'h24: begin
                B_1_round_59[31:24] = SM4_out_12;
            end
            6'h25: begin
                B_1_round_59[23:16] = SM4_out_0;
                B_1_round_59[15:8]  = SM4_out_1;
                B_1_round_59[7:0]   = SM4_out_2;
            end
            default: B_1_round_59 = B_1_round_59;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_60 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_60 = 32'h0;
    end else begin
        BK_0_round_60 = 32'h0;
        case (clk_cnt_all)
            6'h25: begin
                BK_0_round_60[31:24]= SM4_out_3;
                BK_0_round_60[23:16]= SM4_out_4;
                BK_0_round_60[15:8] = SM4_out_5;
                BK_0_round_60[7:0]  = SM4_out_6;
            end
            default: BK_0_round_60 = BK_0_round_60;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_60 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_60 = 32'h0;
    end else begin
        B_0_round_60 = 32'h0;
        case (clk_cnt_all)
            6'h25: begin
                B_0_round_60[31:24] = SM4_out_7;
                B_0_round_60[23:16] = SM4_out_8;
                B_0_round_60[15:8]  = SM4_out_9;
                B_0_round_60[7:0]   = SM4_out_10;
            end
            default: B_0_round_60 = B_0_round_60;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_61 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_61 = 32'h0;
    end else begin
        BK_1_round_61 = 32'h0;
        case (clk_cnt_all)
            6'h25: begin
                BK_1_round_61[31:24]= SM4_out_11;
                BK_1_round_61[23:16]= SM4_out_12;
            end
            6'h26: begin
                BK_1_round_61[15:8] = SM4_out_0;
                BK_1_round_61[7:0]  = SM4_out_1;
            end
            default: BK_1_round_61 = BK_1_round_61;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_61 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_61 = 32'h0;
    end else begin
        B_1_round_61 = 32'h0;
        case (clk_cnt_all)
            6'h26: begin
                B_1_round_61[31:24] = SM4_out_2;
                B_1_round_61[23:16] = SM4_out_3;
                B_1_round_61[15:8]  = SM4_out_4;
                B_1_round_61[7:0]   = SM4_out_5;
            end
            default: B_1_round_61 = B_1_round_61;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_0_round_62 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_0_round_62 = 32'h0;
    end else begin
        BK_0_round_62 = 32'h0;
        case (clk_cnt_all)
            6'h26: begin
                BK_0_round_62[31:24]= SM4_out_6;
                BK_0_round_62[23:16]= SM4_out_7;
                BK_0_round_62[15:8] = SM4_out_8;
                BK_0_round_62[7:0]  = SM4_out_9;
            end
            default: BK_0_round_62 = BK_0_round_62;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_0_round_62 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_0_round_62 = 32'h0;
    end else begin
        B_0_round_62 = 32'h0;
        case (clk_cnt_all)
            6'h26: begin
                B_0_round_62[31:24] = SM4_out_10;
                B_0_round_62[23:16] = SM4_out_11;
                B_0_round_62[15:8]  = SM4_out_12;
            end
            6'h27: begin
                B_0_round_62[7:0]   = SM4_out_0;
            end
            default: B_0_round_62 = B_0_round_62;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        BK_1_round_63 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        BK_1_round_63 = 32'h0;
    end else begin
        BK_1_round_63 = 32'h0;
        case (clk_cnt_all)
            6'h27: begin
                BK_1_round_63[31:24]= SM4_out_1;
                BK_1_round_63[23:16]= SM4_out_2;
                BK_1_round_63[15:8] = SM4_out_3;
                BK_1_round_63[7:0]  = SM4_out_4;
            end
            default: BK_1_round_63 = BK_1_round_63;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        B_1_round_63 = 32'h0;
    end else if (cfg[2:1] == 2'b00 || cfg[2:1] == 2'b01 || cfg[2:1] == 2'b10) begin
        B_1_round_63 = 32'h0;
    end else begin
        B_1_round_63 = 32'h0;
        case (clk_cnt_all)
            6'h27: begin
                B_1_round_63[31:24] = SM4_out_5;
                B_1_round_63[23:16] = SM4_out_6;
                B_1_round_63[15:8]  = SM4_out_7;
                B_1_round_63[7:0]   = SM4_out_8;
            end
            default: B_1_round_63 = B_1_round_63;
        endcase
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_2 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_2 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_2 = sbox_kout_aes_192_clk_2;
        endcase
    end else begin
        sbox_kout_aes_192_clk_2 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_7 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_7 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_7 = sbox_kout_aes_192_clk_7;
        endcase
    end else begin
        sbox_kout_aes_192_clk_7 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_c = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_c = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_c = sbox_kout_aes_192_clk_c;
        endcase
    end else begin
        sbox_kout_aes_192_clk_c = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_11 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_11 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_11 = sbox_kout_aes_192_clk_11;
        endcase
    end else begin
        sbox_kout_aes_192_clk_11 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_16 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_16 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_16 = sbox_kout_aes_192_clk_16;
        endcase
    end else begin
        sbox_kout_aes_192_clk_16 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_1b = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_1b = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_1b = sbox_kout_aes_192_clk_1b;
        endcase
    end else begin
        sbox_kout_aes_192_clk_1b = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_20 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_20 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_20 = sbox_kout_aes_192_clk_20;
        endcase
    end else begin
        sbox_kout_aes_192_clk_20 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_192_clk_25 = 32'h0;
    end else if (cfg[2:1] == 2'b01) begin
        sbox_kout_aes_192_clk_25 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_192_clk_25 = sbox_kout_aes_192_clk_25;
        endcase
    end else begin
        sbox_kout_aes_192_clk_25 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_6 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_6 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_6 = sbox_kout_aes_256_clk_6;
        endcase
    end else begin
        sbox_kout_aes_256_clk_6 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_9 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_9 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_9 = sbox_kout_aes_256_clk_9;
        endcase
    end else begin
        sbox_kout_aes_256_clk_9 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_10 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_10 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_10 = sbox_kout_aes_256_clk_10;
        endcase
    end else begin
        sbox_kout_aes_256_clk_10 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_13 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_13 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_13 = sbox_kout_aes_256_clk_13;
        endcase
    end else begin
        sbox_kout_aes_256_clk_13 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_1a = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_1a = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_1a = sbox_kout_aes_256_clk_1a;
        endcase
    end else begin
        sbox_kout_aes_256_clk_1a = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_1d = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_1d = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_1d = sbox_kout_aes_256_clk_1d;
        endcase
    end else begin
        sbox_kout_aes_256_clk_1d = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_24 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_24 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_24 = sbox_kout_aes_256_clk_24;
        endcase
    end else begin
        sbox_kout_aes_256_clk_24 = 32'h0;
    end
end

always @(*) begin
    if (!rstn) begin
        sbox_kout_aes_256_clk_27 = 32'h0;
    end else if (cfg[2:1] == 2'b10) begin
        sbox_kout_aes_256_clk_27 = 32'h0;
        case (clk_cnt_all)
            default: sbox_kout_aes_256_clk_27 = sbox_kout_aes_256_clk_27;
        endcase
    end else begin
        sbox_kout_aes_256_clk_27 = 32'h0;
    end
end

endmodule
